��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;������Z�������$m|���P�b
��������[b�	��e���}����K�Bs(�����=���m�m�1H�ῗ=�ZiJ�)ڝ��g��ˌa ��@��T�n�ҿYH�Q5r�@��2	��Vn��YŲ�N���,X���\ԥA�&�a��A�2K��s��VZ5���8��ש�4RO���m������&���N�N�B#�$<�����m_lO� �8[S���,�c�/��/���}�;�Aj7Y������3{,k�I�"�r��Y�U��<��M���${�� ՗WNX�J-�%5��aH����S�-!G�e�?�.ή3�pC��}���������Y�;��8�a~�l@ߥ��k�Cv��#���/�҂�&���B�͗Ԯ*Q����P�"��c=�vb�!ф�����$N=�;q����[��$����-Ǹa�WX�s���9:����"�����]f"-�o`�Y]�K� J�xE{�,'����l��;j�m��������q�ex꺑��Ϋ��j7Ţ8��=� ��6�^ڱJ�XF�;��q.�^�ig��܏X`c���<C�g�r�R	�&�ü�C,����\`�Ԛ��U2ڼXQ�l>V&�f۹o��BW�V~ u���c�x����E�Uxd�Tgu���S4��!E��c�L]�c��5�V�i5ցw���g=KH[��z���}���K١�*�Y��`6Nf������&�&$O�GU.>
����x *�胜��T�a�
&�}|M�!QsGD�ݳ��k��<���������/Q�H�努��3|�('F�^J� Xx|V���&�<Y���a�<яL���V�?:�57<�	���o���ec��̫���\��7]Xc�YmK`$?މM �R�.ZD(���θ�:��jH,.���v7?<m-��>NLh��x�:�����S�A,I�]�h�o:QI�z�r��k�C0A6<V	����Ѕ(��R�_�L��}���U�"=�'�2�!~�VT����&��N8ax�Ȑ��I��.�,}!��ig^�p�jӋ� �QǤL�7KU�8fɂH��3�.Ql�+.}��w�I�d��f�DB�5a�ms{}�#�^��X3}1���=k�I�9p�xC�(��w�� ���v�V5EY�w���4�q�5��6��N*�}@�B������"0��Wk]��΄v1�l���	$t��Z���Z�B�P�͜�i���F�T~
�8r*��P�L1����ݬЛ��=!^�� �P6�au��<`�������ڄ�
����qi�'��E1�1\"�È)�����꫞4y2�yh��>�N���3Y����BOu/,O2~4��*�;���o��g��_]-�o�Z��o.G7�*kY�
�P���$`rOVp��E��bd� �Dhv���7^R�.�o��k�g���30�y?b�j�k� u�Sm8YU�>�ؚe�T�\��Q؂��'n����_}}��.+����Z�4k���>�M�U8�%Z��mt����=��0�G����T!�s���V(� ���5g�������������J�z���Ȗ2��4t�����8od,5%[b��(HPɞ-�V7�$�r���oq��֝�%ĺփ �b�0��u�tCi�� u�AԂ���>�ܠ���&�|D�2��i�m�V�!�C*�0��x��Y�q�>�L��g��Qh!r�!_Д��E��灇�1hmA	���>��x�m=p6��7�Vm6�g/C�Ƭfe�������ƹ}��<��Q��k�/B��0��oW����,��g[���{��۸y�qK/�N)ˉm�"�٣��gIH�k�}����ְ��v�H��#�MB�U�z4��2ֻ�]m)�����G��B�hx��-2D�|3*��ǥW�oB��y_ ��KR����8�^��u��:��z�G�;�
ۊ��7����e��VSB��z7����֚�.�BI�Q���f6��S��m�Iq�!����J��.��_�����>8]�(|�������f<2�,�цM8�)�����ǦC�S���d�r��(5��������6�F���<�o�#��0��U6L�<�B3�r��:ǵ�6>�Ӄ�-��͏�w�u'�S�FOr���Q�>W�t��"��R
�4�i��2�W j�~�X�'�\Q0|���!��h�MF�&�$�g�id�	-+�+x5�/�pb`Q0�'�
W�
���N;�I��Y�~�9j���9R�>_�I|�7Zo?��Zz.����������,W�z�,�?1�� ���@���f�d��M�{�9,�
d��=��"��(Q(Fu�M ��cx��i�̋*q��Jw;�g�ȼ_����j��JZ�BF_�v�\y�A����e����N_�3Ԯ�Ñ�����n�
F�>�)�T�QaI^R��k8B$\8S���oHZK8#`8�7�!?�S?��6ij?��Θ*��u��DX]w���+��ˈ����B2뙦����ݱ�N�Gj�{�*�x���3��=^!p_�ّ!}jNȖ�6�o���������Z���	�.��=��K5�C=���9���a�w5g���ov�E�[+~�'�	���R�_[N2�ЪE�}���_z������(W��*�y��%�D{.F�U�۟"\k���w*K�[7�&%g���=qX���߭;d"�ͺ0?G�d�w�J�X�ͯ�����f�S��[��C���n�b�P���?�F�l�S�}�Ռ���8��O�ZjrY]ʔ���f)rѡ;��]��C����	�p6x��SKмֆ��l�{�!�A�\Ʊ��`Sv���	0_NU����SAZC��O@	��|���X���J�L$k;�f��-䅧L�w�Z�Qb���e�%�.�����gQ#��?�����������?Y�\��l�N�	4`�K�EQ���:<ԣ�w�q���&��;��|�4TuMGWK�=Si��t#j�&��c`$�����+��\�ܮ/�6�FD�ӃA��Wp�r�����he,8�I��UN���Q&��T�>m���Α5�7Rֵ?�7��^l ��x��֨T�}����X�W�5mc�r�û{!��.�w2��VD:�y��E��"������҂�X��
T*P����wr�UKIi2����ofq�u��|4�.� Et]l2:�ͣ��ep���i΄��%����E��sJ��8��Nш&cxa1;�G�j	��snj�<o7�R�O��&'ʦ+ͥx5�%��}��4�P���Wu��h�������ץ�b�?�K�U����.�> L�����r�E�2\k$�x�$;��.3�j�馡��MZ��Q[78=.��	�"Mo+Ӿ��6�,�w(�[9�(ae��Trc/��ⴳ��p��do�4�H�WB"�:�o.�����Cj4����ݬ���"�]���r��J+����:��SVU�^$�%�i��yeP�F��S?VbS�>j��(���"�*� ^!Y��xq��:�y*��N���7��Ũ��Q�z����}���)�� ���D6 ��Fʵ�d,��k��[����?eeD�L��P/�/��`M��K�~�������@��*
�n��{�t\~���� c��|����&���bC����e�-� �7��/��V�Z�%"�H�~�꿶��S�Ά�����ݍ�L�����V��#�_
���L�|ea��:�z۾]aXDVWIW�t���@h��}tI�!8�'|Q"���6�/y8NH��"ڃ��4QF�c��,�B��/�0�x���f��!'P�OH�-��0��n�!%��6�pKph|�z��9Z��] �	t�J��R�F@����F���
�:�Kmxe���P��U��~�(Ef/.��T��bt�BPr;��d1�z)M��:r^��c1uǧ���\q2D̓�-�=��&rz�-ˣi�fC�n��l'|�=����D��m(�)Ɉ��fֱJ���7h����f������=o�K��łJ��7W��*�eiJ��>/J�I���o8��M!��^Y�cgز&�O��2泍�mhs����}[ك�ac�""�y=���*���Q�K�����J�5�w��-u���>��{�M���J�KS5 <!<ϸ�����Z�Z�2y�~���?ph�T�����%#-J��+�`ԺЀ+lV�L�H��[�y�5�X�h�7sa�ۼ��2��TFȜ���8:���ծ�϶C��
˅�P[���.�ݶ��q��Lw�p.P^�W;��ȍz��}[���Hln¬%I�"p��g���P��%D-߻�'/�����A�$�0ꏇiVl�q.�q��рw̯�-H��oQ��������l��C��=��c/֍�*X���������!��wЛ�>T~u�-�Ltɸy�"�����s)�E3Si�X�u�zR]4;3d�QD�����%;."gF[ֈq@����J�*:�Q��9���0���x��@�2ց6g���BL4�*��݀�����Fp-���Ij�"����0�kz�Y�弖�'���cu����\a�إ���f;7l	��}�?���?��w����d��$'��5'�1���l�$��d�J����n�j7��P�3MOj����7�Z�$��]���7�▻/h�%tǏ'r��η�yخB��|�62���Voz�r!��gc����H������6N�5��=~�-��-1��gGMv�<�tשuV3`p?f�q��:xT�R���)@�}���E�F[9���{�ᝒ��cl��GHi���V�#�se�n��� ����)�>$���h�����u'��������'~a����ZF6�ӝ �K�S�!T���c���u�y9(�/=ФWQ��]��f���N��v�l��[%L��X���b����X5nspz5��P�Z�n<�E��$W���xx���۾��f���!�dA�Α1�)�gi��痃��+����}W�(�%�	z�F�<f�	T�x�v=<��U�v)�SQV/@�b�_P���Mo�R`L\��^]�ezPgj�6�.j��u~���'*���y�F�)]4\v?:�U��e��K��y�{y�Y�����'�G�X �1e��T�3Z�4��{�-��m�Z�Fg MU����a�=P+��v�pCe
�ܼ�;N`H�i*U��SPzd�$�%
d�\�|�8�Mpx�T=6�ꐮ�EE�@Eٍ�����@w��w�G�C��L/��0� �r��I��a�Ӳ`�g�E]:��˜����IC�O%�B�40��&��D��V�?;N"��|Yt̊g����iE���l�w�d\��ɡt��[*�����)�u4Hg5L��h!F��[��s��1�s�T6�����B�;����8�.�y��їډ�C��h5y:�Ǹ�Q���~t����({�_�h����r-�օ�[hmQ�FO̘�kj�u�؍�O�[E�_%Vr7�Fb|�\���G��ʶ�4��)� l�G�j�������fK��7bϗ��������%"QO���4j�y�m�i�f�>�IM\�]E�b���g6ˍ'�W9�C��4�Q�����������'!)�>�J��й�j;6_����@�*�+���`Po�=�>��ZNDƃ�'��G�el�y����M�E���p�	��3�w���:���Ss0(w8~Ȼ���Ѻ�>(�DSS�lR-�Կ�W���� ��ݳ �i�~��1j���nݭ� ^�;�;+n.}/� i�J���=���lb��#K�MH������h�;&���� ���Ѥ�S�Aeg�����v��A�"�ѓ&�����l���0<?I�{P��.�d������WS�}��&�D�dE��`!�7�~��-e\��Ԡ��6���Lx
�j�UJ��@��J���l�W�U�<��g*϶���p��AdZw=C�����dL��F��r��dm�fE�/�6�D���L�tY����g�I�:ٮb��_��!��y3ڙ�(�M(<���@;�EM[�A	BZ��^|�!V\�d�^2��k�{)�8�@����*a�3�2}=�Y[6�!o�=��&X��������ۦ��e#�7���쎝	¨ � O4x��烣ǣ�J��T-����/ȓ��A�ZA΃=)%7ۭp@Y�R�K����ZhF�եS��mln+��j)f�����gI['��H��"��,ؗZXO���&�t�a$n1�s)'�T*���L"���,���Fa�3�l�0�ZiO~����LHt��#`���U�l�ǵ��Q:W	��LEn�:-��b��q5�E�l����M	_�/c�3z*A:��շ�m����%�i�
&
"�D+Tt6P��v<���k�&�-�񝒝�>�_���H5�Y�����p"���h`/�/�2)�'�e��u[�f]����i�����<�;X���b�0�<R2u}߂�xqer��@��Çv/��茤�+&��.#�tA�Y��B� ��qc�����G����w*HF찆\Š��%��5��m�>�O�P��>Y�=����6Ir"H�m��G��E�΅� ���3��R���:N^Ccn}4�9�S���^�@�"ù��kȁ^^��Ą�Q8@)6S0h�6��h�K����_ߪ%����S3�1��	�N~.�C��M�<wU�"�ݴEK���˪
�Gb�`�Z�՝�|��N��.���^ǀ~2J�$��σ]��}�Rj̀b�F�t�(���PB%ߞ:/�h��"����`^=���j	|����M�N����{����@@�?>�M��0�؉͑�����&K��y�7�)�z[�g���8CM \�Q�]��L�F�7��h�]�&�P|:4%��\�dʢDM��d���1�ViC��F��=���`���HWr�mYv��0K@Y��" ��1�X�a������m]���� zM_��gZR�7�$�P��$o���{p��3���J�98f�\��A���2ؖ�C���1\ԩ��ɡ�)�	�k�O�+7_�x]z������Ԋdn�ΤJ��p��A�uL�����o{���`5��{��A�L�!Og�5x��-�ʫ���]���$/+�W�֙����]��!�@С�Ե׆{b��:|Ymmv�xM�Z@	�i����=�`_�R��*�R2����ɂ�(���r�Ȋ��K��,8p��<3�2&���H���RA-����x�k� jv}��`��5��/�؇5wG]��+���1��?�d�^��z�T��X�Υ�"`'%}�s�'e�1/�$A���ף�3�0�9g���*�܋7�a?�#��h��n�v������쟹w���9�Q  ��j��i��~���2��Q|#!�a��F�l;(m/� ���%oͼ3�_�8�V�q���Ȃ�!��vq�(W$�M@����W���x�hCW~/�P{T�G�2��v�@ѿM������"�b��hƗ��]h�-������;��J߫@��������:}��m�����0�u��� �h�6�������o���Nka>e�6a2�Ӊ9���mu���@6#"��'��2�E!`�Q��X�+:�䝀��8�:i,�v��'����eh;cU	�<���h2��6
m%��1�n���u�f2©�r�+�����RaV-�ks�ә ���D#53��{?H�4��ɿ2�a�	����������t�O_u�O�j!v�0�ZIb��h�����.7�\#��t��-�U,���Xd�	S�<��㖃��R-���M��A�< �n��]t�^�o�Q_���m�&6j�Hs��%-px�ى��h�8�˹��b�)�=���E�� �^��>�0��x��n�D�)�a����_�)k�n7�N�:�/>�iB�X͹U��̑t���U9��\O���U\Yg9�y��J��J&�L<0������J�q��fjѥ	�|{����7�|�:�⤗0,�T!I	����1MA�r0�F���7�8g�ґ�p鸽����u,>��8@�×��Q�h��Wn��8�c��&^q� ����/��&��{j�	�����3eV:`I��YO�
��@����-�B��q��5b="��X�ZVY����!(�j�O=B��	h�==�;9�blkZ�I�}n�.�v\W��6��Q9�8�}�	sф�S�6�8�)T3�0��&s��(�:;z\i������ �HeL�A]Hs�}a@� ���apk��OƘ^�ۤQ	�1&��@��QT��)���WN�>��D%nע�l#���j֕c�~��� ,��Z���2O.-�����{TN�M�U;ߕ��v�VHk�K��}��f_�	����F�ڔ/ʠ�(����x@��˔c���5�S�rY�&� ���]�F^И��3CM�L%X���;���	�������Vf�7REw�n]����hMo$G��K�|��a蛶r=�c�Ja���5��{		;�˂�̪N#؛_��/y�e��کK��n"#~o,2XT���O��`^nh J�����./�.`O���a5��S����ؼ���f�յ5:��k���V��&���u�\�)�6�`І���&�����&��f������Mujf�͐��� �BM_4&�4qm��{�R�g��	RؗU<x�yALS��G��`w:4��vސ|�=Z9dR��"L_��b�A�">LЙi^(�#]�Ϲ�D#�F�X�h��Q�j�'��۶�\AA鹉�rcL��D�o�p�S
 ��!���T�]�7�����}�y��c�5����n�$'iS \����(ߓ ��K�}`�'�����E����w���5�-"�8v��X6�̲d~�d��p���wG1���t`��/�Y�<�.����P��-������.�rvե�W�xES�D����/!S���*��j\κ��E�p$��hN;� 	��Jb�g�Q�˃N��8�R^�lJ�=�ǗQO�6����[�w��K���S�ա�39��~��@ͥ��VRja���G����ߐK�jm4�㟩��`F��bt	W���1S5傤��Le�^���`ӑS��2|7��&�"�cGV��5H�j�皆��
o�NL���*|w{ae�K��ǐ�&422��8m������'b�ZX3ؖ��4֮��+�*S����$��O:�t�'u)�LŻ7�#��t��?�^�����?�.�{��(�O��]F�����|�JuW�/[�lf~r/$����+`RT	�#:��n�kԘ�M�]f 5��>b��{4 ��W���o��drn*�������-��I�0����[��^3��2}�<���X/[�"���[d�֑��WZ�IU�L�rN�W��o��KӒd�rG3:a��2��f�XA�X$k�����h/��<1����WG�6�"%�	�wN���\d���=�i�G�:X��n��5Eds��7:��
�/@ӹײL�kd����U��_��L��2vQ��Q.�Y��>�M���3�M��m>��Ų���`6��}�(�0i�O#.�CvQ7����NјszX۬?����z��r��#��Lv�V�qW;���6w.�����n���60������T��EO�������z��Z�r�Q�E��5ZB��߬tr�q>���mi�%#y��I�0�:�*#c(`�l�>�rm���<���Oh7]~3�(�Ȓ�������y��͠F�,�za�\�fz��z��M��	+u���|�u�Ճ�/��ot�G����'��K/C~xf���*� 1R|�,�jsl�W�&�1,Tj�R#-]���#º��d��rs*.������R;"����(|.�0fV˽��'+��G�_��]���*;���T��=��,��t���Œ��w[���¾^��~�����}M8��m0r�ԄU@�_Dq�l'�����y�c6
ĭ��A��y�(�P��Q�Y}�6�ψ�4BV�4��վ����w<�|����rf�-ж:*(z���&��5)������<@U1Z每���4�C�)���y�:�eD�����#�1��V��y$�S��V��N���bq����_��mE���P��'V�O��`2AY]��,N^&�#=�M9����9���jN��
۹�� �����
j~�P�p��3�L|ڕ���p;:m�Ek��/w����1lv�״}@0o���a{��T��h��>(�?�F�B��$�����M���3��K�9E�U��A����_�z�`4�g�!���Ǭ\�>������Vu'�����e�5�?��]��t�m�u��ts�9����k���*���$jY0�I�!{hD��Ň���]��eo_:Q��a��EU�P����/ǅ\Qp�o<��%6Ƥ�c�N���[N�1w{�]C0#�!����3�Pq
8�Ӟn癋[�K ���=��ls;v��i��DYq�������A$Z���5��`@�R�r'qk�!f ��:�4=�k�'z4Ծ������:F�M�e�왒J�%���������o$�O@�?��C����������4����;�\=�> ��R^ ��F���@'`�X�|S�)�M�9���&��ǐN�2��	��V��F Όg����mб����{c���A��Y�.돣�~��ٓ֝�j1�X��<EVㆌ�sE�f�X����A�Ҕ�V'ǵ�9)�?�n)����;��4ک��y'Sw�	��̸鉓�(p��f��y�w����㓗�d]h��UK:�(K��f��� �J�}��Zc�^�> O9��$��6��}̬��0��✦L���9rY'����A��U"�?�Jp	������M�u<���-�Ij�E�VĤil_㉿:i��VW��i�����Ш�>21g�
�uZ�5�B�CY��8��M#࣒O���0o�`:��`�G�F�c�߼@�H��'}v�����<u-З�{��L;IG�*�����B$l�Kf���4�1�*�����6}>�׭�m�,6�0�DP=+I('E��t�m��h�-o,�L��2���/�@�����%quPZ�B�
���-�K�#$�Nz!�Qf��(ʓ�rYGX����kƈkd�o}�g;?��Uαw�&߽ը�E�꒶�?'o�7,�
�>�F��iOK�Y�_�ڬz�O�`m�T�&H��������y��?Du��v��U���w����m�̣S l鮶��Dc�1���P���Bl}�7[8ݿ��Y4.�[����a�;����&P�ߜ�73�4��t跳=�2�x�x��k&�y��MP�� ��}X�X[z��L�����V����w�=�"�hj8�/͚ω4;`��.o��̿~���0�m�#G7����g��$���&bz��s
vY;�?�8Tq����
$�b�^mA
u�c)�޻L���8?5�u�_�G,�Q���M��K�h�␱�6
��zϟc�yg0�"~���D�j���K�I���5.ɘ.�������}�3���Өu���E�z�Es)��{��:�g��7P��y�â�� �p�7�֔�<�l�����2n��sW�J���97���9�a'^�W|۝�h�l;g{:��E�^q~Y���WF�j�D�m�5뻮&�{��<2I���5K�����|���ԟ?���d28��>���!�N���c�e�ӊ��T^���yF1N���;WŇ]&ce�Q�r�g��ЮL��]�k�p}��e4��Hh@�/]$p�4مb�M]ȡ���v��Gcz�}�����L�t"C>�M�:*t��'��HG�S3BI-W�8v��*�%��]�`��Wա����q��L�O��q���yUe��{�MI|B�*��P��#��1dX�I炤*�G�fx}hy����%��s�G��h�R�Ӣ5�t�k��N05���_�-%}t��W�P��_*�#�!�/��ߤ�<#�x�����6����WM3��%�(�i��ʁ�(��HBw(� ߸�!8~M"���B8��I��o����ǔ���ߪ݁�#|�k+�s?�lW� �~t%���ƨw;�!������-N�>;�n)ܢ��H�1�v��Q3&��G8j�n"D�(�Ƙ�A�(��wE���N��U���Y��pg�S�*|�I��גl8ր�aO�j�
$)$2z�T�u���l��~� �m4��/:2Z��y�%ɥ���a9�� 5"��HEgQ���Ȋ5���ڀ"zz�K�m*EMoÌs��Cq�>�)K�"=�k!��'v8��!i���K��g�6��A�Q���o�'$��[�譪���N�D*]4��	�=7���{�L��Z�����*VQI��0��%�ɋ�d�S�y�=��2�g���0DnP	��hH���aAu஘�LI���)�8�����#�
&	�A<���ѬP"]�3,iΙ���~�X�����5�i�U�B�=�t/Wf*��a��3;yN�X"����$���N�`nv@�!�mS�He+��� �v�����Q�]Ee��Ga��R�_A٠�=i����|\�J�+���zZ�9ԣ;�Q-��V��z�M�\BUc�(�$�ښ��^�a3�)�p9�S�x����/�t���[ַN��%�O=DV�2�!`�*�]�t��=b���K��K4"Ɉ��zΈP�*5��B��p9�3�Ѿ��4.f����O*8�$qs��l��ĕo�q3�ϳ�R�ɟ��p<D5>i���1�ToFJv���H�d��^�t���%н<N��+Zb��;�Px¸[ξ�G���莢�����AZ�)�QA��N�Ox]\��%��AkncnCkf�":5<D#]����Ⱦl8x�f4TZ�Zd���VJ�d���{����gq��z���;�ӱA�H(פ�'39Css:�lJ���q���ժ.��m�����S��1�8��Q8��(����!8���K/O�AAg���*Oz�a4�I;m��xZ��l��!�k�(`s��^�T�������]�����0�d-���A��]�W�~|���uy�Ɯ�e�����*)���ߛ}�����P�.H���ݓk	���r�}�T��v��,ԙi���_�h�ƞP��k�N�I3���@�6��
W�ϳ���_��P���Nv�W�Æp4;�J�O���7�<�M�t}C�_��^��Oe/x5s�X�O�x䋼N�wˏl��!��r�&��6��&j���>�/E	�0�����~�ݐ8=rOԍJ#ˡ�c�z�*�=��;�+�q,��WN�f_5ښHw�Ci��()=5駉B�Ĵ��|����$R}ҹp�w�]9��nБ.�4��N�.���Ú�-]D�L?A�%G�c}��zRIR�T#�ސǬ���V�sθ�:j$�m�:'��{|�?�/ZBfv�����@#`|�L���4Դ���T�����&e���SD��#���u�q���/X	�b4���_3��$�j�0�s���Y�t��VQAs�m��H�8ks�r��2~�=��?�q�ui`?�L9���
��� #'u!`���u互��V�	 �CCg��c閃ͮF2HS�m6fvMT�f5���R�v�Ƹ�o(ˉ��㷇��k
�%J�{�~�(|�^ibh}p�����H2�Ў~S��/{�K�O!=��؏`i��P��J�g�lax:���c�MN����:Y�=7	��D���FP�6�!��"�8����ù �~���R�v�(S�O{(]���3C�
W���Z�"�,��,��'�<�%]tS�l �i�v�8��n��n�����K�F��~D�Xl�������?e*�����ȣ�ָ�2E�OpS�Z7��b���Ң��q<9�)��T7�p�F��jvȐ��x =�ǡ�P��/�p8+*c�ރ��y�K�&JӼUKT��j�^�M_�# �33o��,j�.U���g�?��	ϒ�6��W)��b��Ey�c�t�
�_�y���e:� ��W���� �ʋJ�;�W��� ��h��I���R��u��s3�K�~��wMW���j_	��_n �M���E瑧�1��}A>���G4�-F�q�h�|��<qKTUc��b!��ˆ��kU��_1�,����W�:�����_;�k4�.F��PW��K�q~'b���֤-"`��yp;�쭻�ӂ�\�dz�t:Rdk�:�Z�ֽ
��S��r�D�Q���)�YU=��^޽ ���<��ߙ�n��R�}z��a[>���hX�ce�`&�$�'Ȧ�N�E�\Fٸ��5������ȿ��.�h�$�(;Va����Rޕǎ>�b��W}�����SA���%�lcDts�Ya�^��a��e=��s"�p�`�r-X�C�*�'��%K���!L֞�!�����D��1���=�h���pj��s�kM�c�7G~�n��Y7�Ȼ�5b�0���$���q�v�%P��@��{�̶���҃C��J�PC�g~����)��Y�鴢j.����[���˂+���ꪬ�ױ����c�����֙����7�[j��bS�b���F��[�����0-�.e�E����զRE�F�]�t&�����b&��{��o?��Q�E�U�۩6��VG}irq�oe����d�U�Y�L*u�Hʛ�P�̴C�E6ȣ2�����d1x�d;��tp�&��]z]������R���*]���{Z���U��' '�[�s�7��#�X ��l�ݵ�u�T�b%�y�4��H��ya-] �A[�J�#]T-��ד�w7�奩A�uC���[��_���-��M��4Q��ۛ�R�7xW�]��Mfi�p:�����I1 ��]�^޿{B^�V�d�����