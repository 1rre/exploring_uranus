module EdgeDetect(
  input         clock,
  input         reset,
  input  [10:0] io_x,
  input  [10:0] io_y,
  input  [7:0]  io_px_in_r,
  input  [7:0]  io_px_in_g,
  input  [7:0]  io_px_in_b,
  output [7:0]  io_px_out_r,
  output [7:0]  io_px_out_g,
  output [7:0]  io_px_out_b,
  input         io_line_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] px_buffer_0_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_0_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_1_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_1_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_2_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_2_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_3_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_3_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_4_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_4_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_5_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_5_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_6_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_6_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_7_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_7_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_8_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_8_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_9_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_9_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_10_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_10_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_11_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_11_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_12_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_12_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_13_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_13_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_14_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_14_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_15_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_15_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_16_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_16_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_17_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_17_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_18_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_18_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_19_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_19_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_20_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_20_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_21_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_21_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_22_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_22_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_23_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_23_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_24_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_24_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_25_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_25_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_26_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_26_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_27_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_27_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_28_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_28_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_29_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_29_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_30_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_30_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_31_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_31_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_32_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_32_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_33_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_33_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_34_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_34_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_35_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_35_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_36_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_36_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_37_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_37_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_38_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_38_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_39_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_39_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_40_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_40_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_41_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_41_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_42_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_42_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_43_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_43_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_44_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_44_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_45_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_45_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_46_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_46_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_47_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_47_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_48_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_48_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_49_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_49_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_50_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_50_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_51_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_51_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_52_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_52_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_53_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_53_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_54_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_54_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_55_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_55_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_56_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_56_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_57_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_57_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_58_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_58_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_59_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_59_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_60_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_60_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_61_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_61_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_62_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_62_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_63_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_63_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_64_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_64_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_65_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_65_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_66_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_66_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_67_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_67_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_68_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_68_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_69_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_69_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_70_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_70_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_71_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_71_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_72_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_72_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_73_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_73_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_74_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_74_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_75_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_75_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_76_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_76_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_77_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_77_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_78_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_78_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_79_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_79_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_80_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_80_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_81_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_81_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_82_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_82_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_83_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_83_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_84_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_84_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_85_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_85_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_86_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_86_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_87_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_87_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_88_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_88_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_89_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_89_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_90_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_90_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_91_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_91_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_92_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_92_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_93_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_93_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_94_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_94_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_95_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_95_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_96_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_96_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_97_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_97_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_98_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_98_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_99_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_99_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_100_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_100_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_101_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_101_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_102_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_102_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_103_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_103_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_104_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_104_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_105_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_105_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_106_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_106_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_107_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_107_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_108_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_108_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_109_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_109_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_110_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_110_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_111_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_111_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_112_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_112_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_113_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_113_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_114_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_114_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_115_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_115_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_116_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_116_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_117_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_117_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_118_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_118_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_119_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_119_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_120_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_120_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_121_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_121_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_122_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_122_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_123_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_123_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_124_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_124_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_125_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_125_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_126_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_126_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_127_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_127_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_128_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_128_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_129_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_129_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_130_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_130_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_131_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_131_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_132_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_132_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_133_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_133_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_134_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_134_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_135_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_135_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_136_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_136_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_137_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_137_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_138_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_138_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_139_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_139_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_140_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_140_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_141_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_141_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_142_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_142_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_143_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_143_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_144_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_144_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_145_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_145_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_146_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_146_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_147_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_147_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_148_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_148_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_149_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_149_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_150_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_150_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_151_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_151_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_152_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_152_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_153_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_153_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_154_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_154_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_155_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_155_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_156_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_156_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_157_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_157_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_158_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_158_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_159_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_159_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_160_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_160_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_161_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_161_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_162_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_162_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_163_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_163_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_164_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_164_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_165_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_165_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_166_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_166_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_167_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_167_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_168_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_168_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_169_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_169_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_170_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_170_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_171_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_171_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_172_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_172_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_173_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_173_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_174_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_174_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_175_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_175_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_176_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_176_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_177_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_177_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_178_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_178_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_179_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_179_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_180_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_180_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_181_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_181_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_182_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_182_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_183_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_183_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_184_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_184_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_185_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_185_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_186_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_186_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_187_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_187_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_188_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_188_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_189_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_189_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_190_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_190_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_191_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_191_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_192_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_192_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_193_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_193_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_194_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_194_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_195_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_195_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_196_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_196_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_197_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_197_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_198_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_198_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_199_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_199_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_200_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_200_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_201_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_201_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_202_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_202_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_203_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_203_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_204_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_204_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_205_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_205_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_206_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_206_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_207_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_207_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_208_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_208_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_209_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_209_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_210_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_210_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_211_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_211_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_212_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_212_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_213_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_213_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_214_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_214_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_215_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_215_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_216_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_216_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_217_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_217_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_218_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_218_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_219_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_219_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_220_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_220_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_221_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_221_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_222_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_222_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_223_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_223_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_224_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_224_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_225_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_225_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_226_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_226_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_227_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_227_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_228_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_228_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_229_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_229_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_230_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_230_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_231_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_231_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_232_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_232_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_233_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_233_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_234_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_234_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_235_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_235_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_236_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_236_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_237_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_237_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_238_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_238_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_239_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_239_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_240_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_240_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_241_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_241_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_242_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_242_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_243_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_243_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_244_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_244_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_245_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_245_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_246_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_246_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_247_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_247_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_248_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_248_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_249_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_249_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_250_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_250_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_251_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_251_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_252_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_252_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_253_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_253_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_254_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_254_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_255_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_255_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_256_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_256_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_257_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_257_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_258_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_258_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_259_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_259_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_260_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_260_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_261_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_261_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_262_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_262_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_263_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_263_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_264_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_264_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_265_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_265_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_266_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_266_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_267_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_267_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_268_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_268_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_269_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_269_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_270_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_270_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_271_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_271_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_272_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_272_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_273_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_273_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_274_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_274_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_275_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_275_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_276_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_276_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_277_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_277_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_278_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_278_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_279_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_279_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_280_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_280_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_281_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_281_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_282_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_282_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_283_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_283_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_284_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_284_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_285_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_285_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_286_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_286_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_287_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_287_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_288_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_288_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_289_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_289_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_290_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_290_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_291_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_291_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_292_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_292_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_293_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_293_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_294_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_294_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_295_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_295_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_296_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_296_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_297_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_297_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_298_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_298_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_299_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_299_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_300_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_300_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_301_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_301_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_302_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_302_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_303_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_303_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_304_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_304_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_305_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_305_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_306_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_306_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_307_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_307_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_308_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_308_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_309_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_309_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_310_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_310_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_311_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_311_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_312_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_312_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_313_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_313_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_314_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_314_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_315_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_315_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_316_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_316_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_317_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_317_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_318_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_318_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_319_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_319_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_320_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_320_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_321_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_321_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_322_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_322_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_323_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_323_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_324_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_324_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_325_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_325_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_326_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_326_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_327_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_327_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_328_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_328_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_329_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_329_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_330_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_330_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_331_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_331_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_332_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_332_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_333_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_333_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_334_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_334_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_335_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_335_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_336_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_336_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_337_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_337_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_338_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_338_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_339_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_339_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_340_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_340_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_341_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_341_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_342_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_342_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_343_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_343_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_344_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_344_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_345_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_345_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_346_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_346_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_347_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_347_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_348_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_348_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_349_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_349_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_350_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_350_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_351_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_351_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_352_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_352_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_353_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_353_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_354_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_354_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_355_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_355_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_356_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_356_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_357_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_357_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_358_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_358_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_359_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_359_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_360_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_360_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_361_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_361_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_362_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_362_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_363_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_363_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_364_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_364_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_365_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_365_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_366_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_366_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_367_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_367_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_368_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_368_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_369_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_369_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_370_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_370_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_371_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_371_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_372_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_372_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_373_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_373_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_374_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_374_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_375_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_375_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_376_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_376_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_377_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_377_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_378_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_378_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_379_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_379_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_380_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_380_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_381_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_381_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_382_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_382_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_383_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_383_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_384_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_384_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_385_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_385_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_386_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_386_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_387_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_387_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_388_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_388_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_389_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_389_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_390_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_390_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_391_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_391_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_392_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_392_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_393_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_393_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_394_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_394_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_395_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_395_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_396_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_396_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_397_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_397_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_398_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_398_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_399_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_399_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_400_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_400_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_401_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_401_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_402_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_402_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_403_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_403_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_404_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_404_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_405_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_405_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_406_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_406_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_407_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_407_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_408_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_408_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_409_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_409_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_410_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_410_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_411_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_411_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_412_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_412_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_413_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_413_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_414_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_414_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_415_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_415_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_416_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_416_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_417_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_417_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_418_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_418_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_419_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_419_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_420_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_420_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_421_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_421_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_422_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_422_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_423_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_423_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_424_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_424_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_425_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_425_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_426_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_426_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_427_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_427_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_428_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_428_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_429_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_429_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_430_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_430_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_431_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_431_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_432_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_432_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_433_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_433_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_434_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_434_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_435_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_435_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_436_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_436_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_437_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_437_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_438_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_438_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_439_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_439_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_440_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_440_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_441_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_441_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_442_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_442_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_443_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_443_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_444_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_444_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_445_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_445_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_446_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_446_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_447_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_447_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_448_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_448_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_449_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_449_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_450_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_450_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_451_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_451_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_452_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_452_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_453_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_453_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_454_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_454_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_455_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_455_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_456_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_456_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_457_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_457_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_458_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_458_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_459_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_459_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_460_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_460_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_461_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_461_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_462_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_462_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_463_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_463_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_464_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_464_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_465_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_465_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_466_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_466_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_467_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_467_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_468_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_468_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_469_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_469_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_470_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_470_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_471_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_471_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_472_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_472_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_473_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_473_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_474_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_474_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_475_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_475_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_476_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_476_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_477_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_477_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_478_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_478_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_479_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_479_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_480_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_480_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_481_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_481_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_482_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_482_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_483_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_483_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_484_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_484_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_485_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_485_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_486_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_486_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_487_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_487_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_488_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_488_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_489_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_489_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_490_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_490_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_491_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_491_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_492_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_492_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_493_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_493_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_494_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_494_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_495_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_495_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_496_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_496_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_497_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_497_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_498_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_498_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_499_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_499_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_500_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_500_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_501_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_501_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_502_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_502_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_503_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_503_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_504_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_504_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_505_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_505_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_506_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_506_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_507_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_507_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_508_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_508_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_509_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_509_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_510_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_510_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_511_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_511_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_512_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_512_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_513_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_513_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_514_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_514_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_515_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_515_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_516_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_516_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_517_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_517_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_518_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_518_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_519_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_519_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_520_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_520_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_521_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_521_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_522_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_522_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_523_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_523_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_524_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_524_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_525_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_525_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_526_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_526_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_527_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_527_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_528_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_528_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_529_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_529_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_530_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_530_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_531_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_531_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_532_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_532_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_533_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_533_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_534_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_534_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_535_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_535_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_536_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_536_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_537_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_537_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_538_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_538_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_539_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_539_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_540_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_540_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_541_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_541_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_542_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_542_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_543_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_543_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_544_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_544_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_545_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_545_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_546_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_546_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_547_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_547_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_548_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_548_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_549_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_549_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_550_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_550_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_551_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_551_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_552_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_552_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_553_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_553_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_554_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_554_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_555_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_555_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_556_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_556_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_557_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_557_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_558_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_558_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_559_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_559_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_560_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_560_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_561_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_561_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_562_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_562_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_563_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_563_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_564_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_564_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_565_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_565_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_566_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_566_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_567_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_567_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_568_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_568_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_569_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_569_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_570_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_570_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_571_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_571_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_572_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_572_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_573_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_573_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_574_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_574_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_575_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_575_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_576_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_576_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_577_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_577_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_578_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_578_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_579_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_579_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_580_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_580_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_581_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_581_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_582_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_582_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_583_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_583_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_584_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_584_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_585_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_585_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_586_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_586_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_587_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_587_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_588_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_588_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_589_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_589_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_590_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_590_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_591_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_591_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_592_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_592_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_593_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_593_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_594_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_594_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_595_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_595_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_596_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_596_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_597_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_597_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_598_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_598_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_599_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_599_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_600_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_600_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_601_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_601_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_602_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_602_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_603_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_603_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_604_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_604_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_605_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_605_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_606_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_606_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_607_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_607_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_608_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_608_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_609_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_609_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_610_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_610_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_611_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_611_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_612_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_612_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_613_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_613_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_614_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_614_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_615_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_615_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_616_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_616_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_617_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_617_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_618_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_618_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_619_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_619_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_620_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_620_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_621_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_621_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_622_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_622_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_623_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_623_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_624_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_624_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_625_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_625_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_626_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_626_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_627_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_627_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_628_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_628_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_629_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_629_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_630_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_630_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_631_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_631_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_632_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_632_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_633_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_633_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_634_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_634_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_635_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_635_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_636_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_636_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_637_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_637_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_638_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_638_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_639_r; // @[EdgeDetect.scala 31:26]
  reg [7:0] px_buffer_639_g; // @[EdgeDetect.scala 31:26]
  reg [7:0] last_px_r; // @[EdgeDetect.scala 32:24]
  reg [7:0] last_px_g; // @[EdgeDetect.scala 32:24]
  reg [8:0] REG; // @[EdgeDetect.scala 12:25]
  reg [8:0] REG_1; // @[EdgeDetect.scala 12:25]
  reg [8:0] REG_3; // @[EdgeDetect.scala 12:25]
  reg [8:0] REG_4; // @[EdgeDetect.scala 12:25]
  wire [8:0] _T_3 = 9'sh0 - $signed(REG); // @[EdgeDetect.scala 37:21]
  wire [8:0] _T_5 = $signed(REG) < 9'sh0 ? $signed(_T_3) : $signed(REG); // @[EdgeDetect.scala 37:25]
  wire [7:0] abs_dh_r = _T_5[7:0]; // @[EdgeDetect.scala 37:36]
  wire [8:0] _T_10 = 9'sh0 - $signed(REG_3); // @[EdgeDetect.scala 38:21]
  wire [8:0] _T_12 = $signed(REG_3) < 9'sh0 ? $signed(_T_10) : $signed(REG_3); // @[EdgeDetect.scala 38:25]
  wire [7:0] abs_dv_r = _T_12[7:0]; // @[EdgeDetect.scala 38:36]
  wire [8:0] _T_14 = abs_dh_r + abs_dv_r; // @[EdgeDetect.scala 39:24]
  wire [8:0] _T_21 = 9'sh0 - $signed(REG_1); // @[EdgeDetect.scala 42:21]
  wire [8:0] _T_23 = $signed(REG_1) < 9'sh0 ? $signed(_T_21) : $signed(REG_1); // @[EdgeDetect.scala 42:25]
  wire [7:0] abs_dh_g = _T_23[7:0]; // @[EdgeDetect.scala 42:36]
  wire [8:0] _T_28 = 9'sh0 - $signed(REG_4); // @[EdgeDetect.scala 43:21]
  wire [8:0] _T_30 = $signed(REG_4) < 9'sh0 ? $signed(_T_28) : $signed(REG_4); // @[EdgeDetect.scala 43:25]
  wire [7:0] abs_dv_g = _T_30[7:0]; // @[EdgeDetect.scala 43:36]
  wire [8:0] _T_32 = abs_dh_g + abs_dv_g; // @[EdgeDetect.scala 44:24]
  wire [10:0] _T_54 = io_x - 11'h1; // @[EdgeDetect.scala 54:41]
  wire [7:0] _GEN_1 = 10'h1 == _T_54[9:0] ? px_buffer_1_r : px_buffer_0_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2 = 10'h2 == _T_54[9:0] ? px_buffer_2_r : _GEN_1; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3 = 10'h3 == _T_54[9:0] ? px_buffer_3_r : _GEN_2; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4 = 10'h4 == _T_54[9:0] ? px_buffer_4_r : _GEN_3; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5 = 10'h5 == _T_54[9:0] ? px_buffer_5_r : _GEN_4; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6 = 10'h6 == _T_54[9:0] ? px_buffer_6_r : _GEN_5; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7 = 10'h7 == _T_54[9:0] ? px_buffer_7_r : _GEN_6; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8 = 10'h8 == _T_54[9:0] ? px_buffer_8_r : _GEN_7; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9 = 10'h9 == _T_54[9:0] ? px_buffer_9_r : _GEN_8; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10 = 10'ha == _T_54[9:0] ? px_buffer_10_r : _GEN_9; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11 = 10'hb == _T_54[9:0] ? px_buffer_11_r : _GEN_10; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12 = 10'hc == _T_54[9:0] ? px_buffer_12_r : _GEN_11; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_13 = 10'hd == _T_54[9:0] ? px_buffer_13_r : _GEN_12; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_14 = 10'he == _T_54[9:0] ? px_buffer_14_r : _GEN_13; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_15 = 10'hf == _T_54[9:0] ? px_buffer_15_r : _GEN_14; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_16 = 10'h10 == _T_54[9:0] ? px_buffer_16_r : _GEN_15; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_17 = 10'h11 == _T_54[9:0] ? px_buffer_17_r : _GEN_16; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_18 = 10'h12 == _T_54[9:0] ? px_buffer_18_r : _GEN_17; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_19 = 10'h13 == _T_54[9:0] ? px_buffer_19_r : _GEN_18; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_20 = 10'h14 == _T_54[9:0] ? px_buffer_20_r : _GEN_19; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_21 = 10'h15 == _T_54[9:0] ? px_buffer_21_r : _GEN_20; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_22 = 10'h16 == _T_54[9:0] ? px_buffer_22_r : _GEN_21; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_23 = 10'h17 == _T_54[9:0] ? px_buffer_23_r : _GEN_22; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_24 = 10'h18 == _T_54[9:0] ? px_buffer_24_r : _GEN_23; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_25 = 10'h19 == _T_54[9:0] ? px_buffer_25_r : _GEN_24; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_26 = 10'h1a == _T_54[9:0] ? px_buffer_26_r : _GEN_25; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_27 = 10'h1b == _T_54[9:0] ? px_buffer_27_r : _GEN_26; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_28 = 10'h1c == _T_54[9:0] ? px_buffer_28_r : _GEN_27; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_29 = 10'h1d == _T_54[9:0] ? px_buffer_29_r : _GEN_28; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_30 = 10'h1e == _T_54[9:0] ? px_buffer_30_r : _GEN_29; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_31 = 10'h1f == _T_54[9:0] ? px_buffer_31_r : _GEN_30; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_32 = 10'h20 == _T_54[9:0] ? px_buffer_32_r : _GEN_31; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_33 = 10'h21 == _T_54[9:0] ? px_buffer_33_r : _GEN_32; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_34 = 10'h22 == _T_54[9:0] ? px_buffer_34_r : _GEN_33; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_35 = 10'h23 == _T_54[9:0] ? px_buffer_35_r : _GEN_34; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_36 = 10'h24 == _T_54[9:0] ? px_buffer_36_r : _GEN_35; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_37 = 10'h25 == _T_54[9:0] ? px_buffer_37_r : _GEN_36; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_38 = 10'h26 == _T_54[9:0] ? px_buffer_38_r : _GEN_37; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_39 = 10'h27 == _T_54[9:0] ? px_buffer_39_r : _GEN_38; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_40 = 10'h28 == _T_54[9:0] ? px_buffer_40_r : _GEN_39; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_41 = 10'h29 == _T_54[9:0] ? px_buffer_41_r : _GEN_40; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_42 = 10'h2a == _T_54[9:0] ? px_buffer_42_r : _GEN_41; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_43 = 10'h2b == _T_54[9:0] ? px_buffer_43_r : _GEN_42; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_44 = 10'h2c == _T_54[9:0] ? px_buffer_44_r : _GEN_43; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_45 = 10'h2d == _T_54[9:0] ? px_buffer_45_r : _GEN_44; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_46 = 10'h2e == _T_54[9:0] ? px_buffer_46_r : _GEN_45; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_47 = 10'h2f == _T_54[9:0] ? px_buffer_47_r : _GEN_46; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_48 = 10'h30 == _T_54[9:0] ? px_buffer_48_r : _GEN_47; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_49 = 10'h31 == _T_54[9:0] ? px_buffer_49_r : _GEN_48; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_50 = 10'h32 == _T_54[9:0] ? px_buffer_50_r : _GEN_49; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_51 = 10'h33 == _T_54[9:0] ? px_buffer_51_r : _GEN_50; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_52 = 10'h34 == _T_54[9:0] ? px_buffer_52_r : _GEN_51; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_53 = 10'h35 == _T_54[9:0] ? px_buffer_53_r : _GEN_52; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_54 = 10'h36 == _T_54[9:0] ? px_buffer_54_r : _GEN_53; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_55 = 10'h37 == _T_54[9:0] ? px_buffer_55_r : _GEN_54; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_56 = 10'h38 == _T_54[9:0] ? px_buffer_56_r : _GEN_55; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_57 = 10'h39 == _T_54[9:0] ? px_buffer_57_r : _GEN_56; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_58 = 10'h3a == _T_54[9:0] ? px_buffer_58_r : _GEN_57; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_59 = 10'h3b == _T_54[9:0] ? px_buffer_59_r : _GEN_58; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_60 = 10'h3c == _T_54[9:0] ? px_buffer_60_r : _GEN_59; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_61 = 10'h3d == _T_54[9:0] ? px_buffer_61_r : _GEN_60; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_62 = 10'h3e == _T_54[9:0] ? px_buffer_62_r : _GEN_61; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_63 = 10'h3f == _T_54[9:0] ? px_buffer_63_r : _GEN_62; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_64 = 10'h40 == _T_54[9:0] ? px_buffer_64_r : _GEN_63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_65 = 10'h41 == _T_54[9:0] ? px_buffer_65_r : _GEN_64; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_66 = 10'h42 == _T_54[9:0] ? px_buffer_66_r : _GEN_65; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_67 = 10'h43 == _T_54[9:0] ? px_buffer_67_r : _GEN_66; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_68 = 10'h44 == _T_54[9:0] ? px_buffer_68_r : _GEN_67; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_69 = 10'h45 == _T_54[9:0] ? px_buffer_69_r : _GEN_68; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_70 = 10'h46 == _T_54[9:0] ? px_buffer_70_r : _GEN_69; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_71 = 10'h47 == _T_54[9:0] ? px_buffer_71_r : _GEN_70; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_72 = 10'h48 == _T_54[9:0] ? px_buffer_72_r : _GEN_71; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_73 = 10'h49 == _T_54[9:0] ? px_buffer_73_r : _GEN_72; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_74 = 10'h4a == _T_54[9:0] ? px_buffer_74_r : _GEN_73; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_75 = 10'h4b == _T_54[9:0] ? px_buffer_75_r : _GEN_74; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_76 = 10'h4c == _T_54[9:0] ? px_buffer_76_r : _GEN_75; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_77 = 10'h4d == _T_54[9:0] ? px_buffer_77_r : _GEN_76; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_78 = 10'h4e == _T_54[9:0] ? px_buffer_78_r : _GEN_77; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_79 = 10'h4f == _T_54[9:0] ? px_buffer_79_r : _GEN_78; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_80 = 10'h50 == _T_54[9:0] ? px_buffer_80_r : _GEN_79; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_81 = 10'h51 == _T_54[9:0] ? px_buffer_81_r : _GEN_80; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_82 = 10'h52 == _T_54[9:0] ? px_buffer_82_r : _GEN_81; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_83 = 10'h53 == _T_54[9:0] ? px_buffer_83_r : _GEN_82; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_84 = 10'h54 == _T_54[9:0] ? px_buffer_84_r : _GEN_83; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_85 = 10'h55 == _T_54[9:0] ? px_buffer_85_r : _GEN_84; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_86 = 10'h56 == _T_54[9:0] ? px_buffer_86_r : _GEN_85; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_87 = 10'h57 == _T_54[9:0] ? px_buffer_87_r : _GEN_86; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_88 = 10'h58 == _T_54[9:0] ? px_buffer_88_r : _GEN_87; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_89 = 10'h59 == _T_54[9:0] ? px_buffer_89_r : _GEN_88; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_90 = 10'h5a == _T_54[9:0] ? px_buffer_90_r : _GEN_89; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_91 = 10'h5b == _T_54[9:0] ? px_buffer_91_r : _GEN_90; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_92 = 10'h5c == _T_54[9:0] ? px_buffer_92_r : _GEN_91; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_93 = 10'h5d == _T_54[9:0] ? px_buffer_93_r : _GEN_92; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_94 = 10'h5e == _T_54[9:0] ? px_buffer_94_r : _GEN_93; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_95 = 10'h5f == _T_54[9:0] ? px_buffer_95_r : _GEN_94; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_96 = 10'h60 == _T_54[9:0] ? px_buffer_96_r : _GEN_95; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_97 = 10'h61 == _T_54[9:0] ? px_buffer_97_r : _GEN_96; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_98 = 10'h62 == _T_54[9:0] ? px_buffer_98_r : _GEN_97; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_99 = 10'h63 == _T_54[9:0] ? px_buffer_99_r : _GEN_98; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_100 = 10'h64 == _T_54[9:0] ? px_buffer_100_r : _GEN_99; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_101 = 10'h65 == _T_54[9:0] ? px_buffer_101_r : _GEN_100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_102 = 10'h66 == _T_54[9:0] ? px_buffer_102_r : _GEN_101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_103 = 10'h67 == _T_54[9:0] ? px_buffer_103_r : _GEN_102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_104 = 10'h68 == _T_54[9:0] ? px_buffer_104_r : _GEN_103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_105 = 10'h69 == _T_54[9:0] ? px_buffer_105_r : _GEN_104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_106 = 10'h6a == _T_54[9:0] ? px_buffer_106_r : _GEN_105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_107 = 10'h6b == _T_54[9:0] ? px_buffer_107_r : _GEN_106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_108 = 10'h6c == _T_54[9:0] ? px_buffer_108_r : _GEN_107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_109 = 10'h6d == _T_54[9:0] ? px_buffer_109_r : _GEN_108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_110 = 10'h6e == _T_54[9:0] ? px_buffer_110_r : _GEN_109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_111 = 10'h6f == _T_54[9:0] ? px_buffer_111_r : _GEN_110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_112 = 10'h70 == _T_54[9:0] ? px_buffer_112_r : _GEN_111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_113 = 10'h71 == _T_54[9:0] ? px_buffer_113_r : _GEN_112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_114 = 10'h72 == _T_54[9:0] ? px_buffer_114_r : _GEN_113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_115 = 10'h73 == _T_54[9:0] ? px_buffer_115_r : _GEN_114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_116 = 10'h74 == _T_54[9:0] ? px_buffer_116_r : _GEN_115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_117 = 10'h75 == _T_54[9:0] ? px_buffer_117_r : _GEN_116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_118 = 10'h76 == _T_54[9:0] ? px_buffer_118_r : _GEN_117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_119 = 10'h77 == _T_54[9:0] ? px_buffer_119_r : _GEN_118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_120 = 10'h78 == _T_54[9:0] ? px_buffer_120_r : _GEN_119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_121 = 10'h79 == _T_54[9:0] ? px_buffer_121_r : _GEN_120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_122 = 10'h7a == _T_54[9:0] ? px_buffer_122_r : _GEN_121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_123 = 10'h7b == _T_54[9:0] ? px_buffer_123_r : _GEN_122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_124 = 10'h7c == _T_54[9:0] ? px_buffer_124_r : _GEN_123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_125 = 10'h7d == _T_54[9:0] ? px_buffer_125_r : _GEN_124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_126 = 10'h7e == _T_54[9:0] ? px_buffer_126_r : _GEN_125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_127 = 10'h7f == _T_54[9:0] ? px_buffer_127_r : _GEN_126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_128 = 10'h80 == _T_54[9:0] ? px_buffer_128_r : _GEN_127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_129 = 10'h81 == _T_54[9:0] ? px_buffer_129_r : _GEN_128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_130 = 10'h82 == _T_54[9:0] ? px_buffer_130_r : _GEN_129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_131 = 10'h83 == _T_54[9:0] ? px_buffer_131_r : _GEN_130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_132 = 10'h84 == _T_54[9:0] ? px_buffer_132_r : _GEN_131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_133 = 10'h85 == _T_54[9:0] ? px_buffer_133_r : _GEN_132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_134 = 10'h86 == _T_54[9:0] ? px_buffer_134_r : _GEN_133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_135 = 10'h87 == _T_54[9:0] ? px_buffer_135_r : _GEN_134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_136 = 10'h88 == _T_54[9:0] ? px_buffer_136_r : _GEN_135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_137 = 10'h89 == _T_54[9:0] ? px_buffer_137_r : _GEN_136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_138 = 10'h8a == _T_54[9:0] ? px_buffer_138_r : _GEN_137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_139 = 10'h8b == _T_54[9:0] ? px_buffer_139_r : _GEN_138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_140 = 10'h8c == _T_54[9:0] ? px_buffer_140_r : _GEN_139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_141 = 10'h8d == _T_54[9:0] ? px_buffer_141_r : _GEN_140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_142 = 10'h8e == _T_54[9:0] ? px_buffer_142_r : _GEN_141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_143 = 10'h8f == _T_54[9:0] ? px_buffer_143_r : _GEN_142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_144 = 10'h90 == _T_54[9:0] ? px_buffer_144_r : _GEN_143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_145 = 10'h91 == _T_54[9:0] ? px_buffer_145_r : _GEN_144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_146 = 10'h92 == _T_54[9:0] ? px_buffer_146_r : _GEN_145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_147 = 10'h93 == _T_54[9:0] ? px_buffer_147_r : _GEN_146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_148 = 10'h94 == _T_54[9:0] ? px_buffer_148_r : _GEN_147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_149 = 10'h95 == _T_54[9:0] ? px_buffer_149_r : _GEN_148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_150 = 10'h96 == _T_54[9:0] ? px_buffer_150_r : _GEN_149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_151 = 10'h97 == _T_54[9:0] ? px_buffer_151_r : _GEN_150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_152 = 10'h98 == _T_54[9:0] ? px_buffer_152_r : _GEN_151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_153 = 10'h99 == _T_54[9:0] ? px_buffer_153_r : _GEN_152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_154 = 10'h9a == _T_54[9:0] ? px_buffer_154_r : _GEN_153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_155 = 10'h9b == _T_54[9:0] ? px_buffer_155_r : _GEN_154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_156 = 10'h9c == _T_54[9:0] ? px_buffer_156_r : _GEN_155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_157 = 10'h9d == _T_54[9:0] ? px_buffer_157_r : _GEN_156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_158 = 10'h9e == _T_54[9:0] ? px_buffer_158_r : _GEN_157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_159 = 10'h9f == _T_54[9:0] ? px_buffer_159_r : _GEN_158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_160 = 10'ha0 == _T_54[9:0] ? px_buffer_160_r : _GEN_159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_161 = 10'ha1 == _T_54[9:0] ? px_buffer_161_r : _GEN_160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_162 = 10'ha2 == _T_54[9:0] ? px_buffer_162_r : _GEN_161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_163 = 10'ha3 == _T_54[9:0] ? px_buffer_163_r : _GEN_162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_164 = 10'ha4 == _T_54[9:0] ? px_buffer_164_r : _GEN_163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_165 = 10'ha5 == _T_54[9:0] ? px_buffer_165_r : _GEN_164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_166 = 10'ha6 == _T_54[9:0] ? px_buffer_166_r : _GEN_165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_167 = 10'ha7 == _T_54[9:0] ? px_buffer_167_r : _GEN_166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_168 = 10'ha8 == _T_54[9:0] ? px_buffer_168_r : _GEN_167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_169 = 10'ha9 == _T_54[9:0] ? px_buffer_169_r : _GEN_168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_170 = 10'haa == _T_54[9:0] ? px_buffer_170_r : _GEN_169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_171 = 10'hab == _T_54[9:0] ? px_buffer_171_r : _GEN_170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_172 = 10'hac == _T_54[9:0] ? px_buffer_172_r : _GEN_171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_173 = 10'had == _T_54[9:0] ? px_buffer_173_r : _GEN_172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_174 = 10'hae == _T_54[9:0] ? px_buffer_174_r : _GEN_173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_175 = 10'haf == _T_54[9:0] ? px_buffer_175_r : _GEN_174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_176 = 10'hb0 == _T_54[9:0] ? px_buffer_176_r : _GEN_175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_177 = 10'hb1 == _T_54[9:0] ? px_buffer_177_r : _GEN_176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_178 = 10'hb2 == _T_54[9:0] ? px_buffer_178_r : _GEN_177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_179 = 10'hb3 == _T_54[9:0] ? px_buffer_179_r : _GEN_178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_180 = 10'hb4 == _T_54[9:0] ? px_buffer_180_r : _GEN_179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_181 = 10'hb5 == _T_54[9:0] ? px_buffer_181_r : _GEN_180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_182 = 10'hb6 == _T_54[9:0] ? px_buffer_182_r : _GEN_181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_183 = 10'hb7 == _T_54[9:0] ? px_buffer_183_r : _GEN_182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_184 = 10'hb8 == _T_54[9:0] ? px_buffer_184_r : _GEN_183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_185 = 10'hb9 == _T_54[9:0] ? px_buffer_185_r : _GEN_184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_186 = 10'hba == _T_54[9:0] ? px_buffer_186_r : _GEN_185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_187 = 10'hbb == _T_54[9:0] ? px_buffer_187_r : _GEN_186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_188 = 10'hbc == _T_54[9:0] ? px_buffer_188_r : _GEN_187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_189 = 10'hbd == _T_54[9:0] ? px_buffer_189_r : _GEN_188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_190 = 10'hbe == _T_54[9:0] ? px_buffer_190_r : _GEN_189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_191 = 10'hbf == _T_54[9:0] ? px_buffer_191_r : _GEN_190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_192 = 10'hc0 == _T_54[9:0] ? px_buffer_192_r : _GEN_191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_193 = 10'hc1 == _T_54[9:0] ? px_buffer_193_r : _GEN_192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_194 = 10'hc2 == _T_54[9:0] ? px_buffer_194_r : _GEN_193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_195 = 10'hc3 == _T_54[9:0] ? px_buffer_195_r : _GEN_194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_196 = 10'hc4 == _T_54[9:0] ? px_buffer_196_r : _GEN_195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_197 = 10'hc5 == _T_54[9:0] ? px_buffer_197_r : _GEN_196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_198 = 10'hc6 == _T_54[9:0] ? px_buffer_198_r : _GEN_197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_199 = 10'hc7 == _T_54[9:0] ? px_buffer_199_r : _GEN_198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_200 = 10'hc8 == _T_54[9:0] ? px_buffer_200_r : _GEN_199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_201 = 10'hc9 == _T_54[9:0] ? px_buffer_201_r : _GEN_200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_202 = 10'hca == _T_54[9:0] ? px_buffer_202_r : _GEN_201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_203 = 10'hcb == _T_54[9:0] ? px_buffer_203_r : _GEN_202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_204 = 10'hcc == _T_54[9:0] ? px_buffer_204_r : _GEN_203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_205 = 10'hcd == _T_54[9:0] ? px_buffer_205_r : _GEN_204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_206 = 10'hce == _T_54[9:0] ? px_buffer_206_r : _GEN_205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_207 = 10'hcf == _T_54[9:0] ? px_buffer_207_r : _GEN_206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_208 = 10'hd0 == _T_54[9:0] ? px_buffer_208_r : _GEN_207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_209 = 10'hd1 == _T_54[9:0] ? px_buffer_209_r : _GEN_208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_210 = 10'hd2 == _T_54[9:0] ? px_buffer_210_r : _GEN_209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_211 = 10'hd3 == _T_54[9:0] ? px_buffer_211_r : _GEN_210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_212 = 10'hd4 == _T_54[9:0] ? px_buffer_212_r : _GEN_211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_213 = 10'hd5 == _T_54[9:0] ? px_buffer_213_r : _GEN_212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_214 = 10'hd6 == _T_54[9:0] ? px_buffer_214_r : _GEN_213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_215 = 10'hd7 == _T_54[9:0] ? px_buffer_215_r : _GEN_214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_216 = 10'hd8 == _T_54[9:0] ? px_buffer_216_r : _GEN_215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_217 = 10'hd9 == _T_54[9:0] ? px_buffer_217_r : _GEN_216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_218 = 10'hda == _T_54[9:0] ? px_buffer_218_r : _GEN_217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_219 = 10'hdb == _T_54[9:0] ? px_buffer_219_r : _GEN_218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_220 = 10'hdc == _T_54[9:0] ? px_buffer_220_r : _GEN_219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_221 = 10'hdd == _T_54[9:0] ? px_buffer_221_r : _GEN_220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_222 = 10'hde == _T_54[9:0] ? px_buffer_222_r : _GEN_221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_223 = 10'hdf == _T_54[9:0] ? px_buffer_223_r : _GEN_222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_224 = 10'he0 == _T_54[9:0] ? px_buffer_224_r : _GEN_223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_225 = 10'he1 == _T_54[9:0] ? px_buffer_225_r : _GEN_224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_226 = 10'he2 == _T_54[9:0] ? px_buffer_226_r : _GEN_225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_227 = 10'he3 == _T_54[9:0] ? px_buffer_227_r : _GEN_226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_228 = 10'he4 == _T_54[9:0] ? px_buffer_228_r : _GEN_227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_229 = 10'he5 == _T_54[9:0] ? px_buffer_229_r : _GEN_228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_230 = 10'he6 == _T_54[9:0] ? px_buffer_230_r : _GEN_229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_231 = 10'he7 == _T_54[9:0] ? px_buffer_231_r : _GEN_230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_232 = 10'he8 == _T_54[9:0] ? px_buffer_232_r : _GEN_231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_233 = 10'he9 == _T_54[9:0] ? px_buffer_233_r : _GEN_232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_234 = 10'hea == _T_54[9:0] ? px_buffer_234_r : _GEN_233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_235 = 10'heb == _T_54[9:0] ? px_buffer_235_r : _GEN_234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_236 = 10'hec == _T_54[9:0] ? px_buffer_236_r : _GEN_235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_237 = 10'hed == _T_54[9:0] ? px_buffer_237_r : _GEN_236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_238 = 10'hee == _T_54[9:0] ? px_buffer_238_r : _GEN_237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_239 = 10'hef == _T_54[9:0] ? px_buffer_239_r : _GEN_238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_240 = 10'hf0 == _T_54[9:0] ? px_buffer_240_r : _GEN_239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_241 = 10'hf1 == _T_54[9:0] ? px_buffer_241_r : _GEN_240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_242 = 10'hf2 == _T_54[9:0] ? px_buffer_242_r : _GEN_241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_243 = 10'hf3 == _T_54[9:0] ? px_buffer_243_r : _GEN_242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_244 = 10'hf4 == _T_54[9:0] ? px_buffer_244_r : _GEN_243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_245 = 10'hf5 == _T_54[9:0] ? px_buffer_245_r : _GEN_244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_246 = 10'hf6 == _T_54[9:0] ? px_buffer_246_r : _GEN_245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_247 = 10'hf7 == _T_54[9:0] ? px_buffer_247_r : _GEN_246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_248 = 10'hf8 == _T_54[9:0] ? px_buffer_248_r : _GEN_247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_249 = 10'hf9 == _T_54[9:0] ? px_buffer_249_r : _GEN_248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_250 = 10'hfa == _T_54[9:0] ? px_buffer_250_r : _GEN_249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_251 = 10'hfb == _T_54[9:0] ? px_buffer_251_r : _GEN_250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_252 = 10'hfc == _T_54[9:0] ? px_buffer_252_r : _GEN_251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_253 = 10'hfd == _T_54[9:0] ? px_buffer_253_r : _GEN_252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_254 = 10'hfe == _T_54[9:0] ? px_buffer_254_r : _GEN_253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_255 = 10'hff == _T_54[9:0] ? px_buffer_255_r : _GEN_254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_256 = 10'h100 == _T_54[9:0] ? px_buffer_256_r : _GEN_255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_257 = 10'h101 == _T_54[9:0] ? px_buffer_257_r : _GEN_256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_258 = 10'h102 == _T_54[9:0] ? px_buffer_258_r : _GEN_257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_259 = 10'h103 == _T_54[9:0] ? px_buffer_259_r : _GEN_258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_260 = 10'h104 == _T_54[9:0] ? px_buffer_260_r : _GEN_259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_261 = 10'h105 == _T_54[9:0] ? px_buffer_261_r : _GEN_260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_262 = 10'h106 == _T_54[9:0] ? px_buffer_262_r : _GEN_261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_263 = 10'h107 == _T_54[9:0] ? px_buffer_263_r : _GEN_262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_264 = 10'h108 == _T_54[9:0] ? px_buffer_264_r : _GEN_263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_265 = 10'h109 == _T_54[9:0] ? px_buffer_265_r : _GEN_264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_266 = 10'h10a == _T_54[9:0] ? px_buffer_266_r : _GEN_265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_267 = 10'h10b == _T_54[9:0] ? px_buffer_267_r : _GEN_266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_268 = 10'h10c == _T_54[9:0] ? px_buffer_268_r : _GEN_267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_269 = 10'h10d == _T_54[9:0] ? px_buffer_269_r : _GEN_268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_270 = 10'h10e == _T_54[9:0] ? px_buffer_270_r : _GEN_269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_271 = 10'h10f == _T_54[9:0] ? px_buffer_271_r : _GEN_270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_272 = 10'h110 == _T_54[9:0] ? px_buffer_272_r : _GEN_271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_273 = 10'h111 == _T_54[9:0] ? px_buffer_273_r : _GEN_272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_274 = 10'h112 == _T_54[9:0] ? px_buffer_274_r : _GEN_273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_275 = 10'h113 == _T_54[9:0] ? px_buffer_275_r : _GEN_274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_276 = 10'h114 == _T_54[9:0] ? px_buffer_276_r : _GEN_275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_277 = 10'h115 == _T_54[9:0] ? px_buffer_277_r : _GEN_276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_278 = 10'h116 == _T_54[9:0] ? px_buffer_278_r : _GEN_277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_279 = 10'h117 == _T_54[9:0] ? px_buffer_279_r : _GEN_278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_280 = 10'h118 == _T_54[9:0] ? px_buffer_280_r : _GEN_279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_281 = 10'h119 == _T_54[9:0] ? px_buffer_281_r : _GEN_280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_282 = 10'h11a == _T_54[9:0] ? px_buffer_282_r : _GEN_281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_283 = 10'h11b == _T_54[9:0] ? px_buffer_283_r : _GEN_282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_284 = 10'h11c == _T_54[9:0] ? px_buffer_284_r : _GEN_283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_285 = 10'h11d == _T_54[9:0] ? px_buffer_285_r : _GEN_284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_286 = 10'h11e == _T_54[9:0] ? px_buffer_286_r : _GEN_285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_287 = 10'h11f == _T_54[9:0] ? px_buffer_287_r : _GEN_286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_288 = 10'h120 == _T_54[9:0] ? px_buffer_288_r : _GEN_287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_289 = 10'h121 == _T_54[9:0] ? px_buffer_289_r : _GEN_288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_290 = 10'h122 == _T_54[9:0] ? px_buffer_290_r : _GEN_289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_291 = 10'h123 == _T_54[9:0] ? px_buffer_291_r : _GEN_290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_292 = 10'h124 == _T_54[9:0] ? px_buffer_292_r : _GEN_291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_293 = 10'h125 == _T_54[9:0] ? px_buffer_293_r : _GEN_292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_294 = 10'h126 == _T_54[9:0] ? px_buffer_294_r : _GEN_293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_295 = 10'h127 == _T_54[9:0] ? px_buffer_295_r : _GEN_294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_296 = 10'h128 == _T_54[9:0] ? px_buffer_296_r : _GEN_295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_297 = 10'h129 == _T_54[9:0] ? px_buffer_297_r : _GEN_296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_298 = 10'h12a == _T_54[9:0] ? px_buffer_298_r : _GEN_297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_299 = 10'h12b == _T_54[9:0] ? px_buffer_299_r : _GEN_298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_300 = 10'h12c == _T_54[9:0] ? px_buffer_300_r : _GEN_299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_301 = 10'h12d == _T_54[9:0] ? px_buffer_301_r : _GEN_300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_302 = 10'h12e == _T_54[9:0] ? px_buffer_302_r : _GEN_301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_303 = 10'h12f == _T_54[9:0] ? px_buffer_303_r : _GEN_302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_304 = 10'h130 == _T_54[9:0] ? px_buffer_304_r : _GEN_303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_305 = 10'h131 == _T_54[9:0] ? px_buffer_305_r : _GEN_304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_306 = 10'h132 == _T_54[9:0] ? px_buffer_306_r : _GEN_305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_307 = 10'h133 == _T_54[9:0] ? px_buffer_307_r : _GEN_306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_308 = 10'h134 == _T_54[9:0] ? px_buffer_308_r : _GEN_307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_309 = 10'h135 == _T_54[9:0] ? px_buffer_309_r : _GEN_308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_310 = 10'h136 == _T_54[9:0] ? px_buffer_310_r : _GEN_309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_311 = 10'h137 == _T_54[9:0] ? px_buffer_311_r : _GEN_310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_312 = 10'h138 == _T_54[9:0] ? px_buffer_312_r : _GEN_311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_313 = 10'h139 == _T_54[9:0] ? px_buffer_313_r : _GEN_312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_314 = 10'h13a == _T_54[9:0] ? px_buffer_314_r : _GEN_313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_315 = 10'h13b == _T_54[9:0] ? px_buffer_315_r : _GEN_314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_316 = 10'h13c == _T_54[9:0] ? px_buffer_316_r : _GEN_315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_317 = 10'h13d == _T_54[9:0] ? px_buffer_317_r : _GEN_316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_318 = 10'h13e == _T_54[9:0] ? px_buffer_318_r : _GEN_317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_319 = 10'h13f == _T_54[9:0] ? px_buffer_319_r : _GEN_318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_320 = 10'h140 == _T_54[9:0] ? px_buffer_320_r : _GEN_319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_321 = 10'h141 == _T_54[9:0] ? px_buffer_321_r : _GEN_320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_322 = 10'h142 == _T_54[9:0] ? px_buffer_322_r : _GEN_321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_323 = 10'h143 == _T_54[9:0] ? px_buffer_323_r : _GEN_322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_324 = 10'h144 == _T_54[9:0] ? px_buffer_324_r : _GEN_323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_325 = 10'h145 == _T_54[9:0] ? px_buffer_325_r : _GEN_324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_326 = 10'h146 == _T_54[9:0] ? px_buffer_326_r : _GEN_325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_327 = 10'h147 == _T_54[9:0] ? px_buffer_327_r : _GEN_326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_328 = 10'h148 == _T_54[9:0] ? px_buffer_328_r : _GEN_327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_329 = 10'h149 == _T_54[9:0] ? px_buffer_329_r : _GEN_328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_330 = 10'h14a == _T_54[9:0] ? px_buffer_330_r : _GEN_329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_331 = 10'h14b == _T_54[9:0] ? px_buffer_331_r : _GEN_330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_332 = 10'h14c == _T_54[9:0] ? px_buffer_332_r : _GEN_331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_333 = 10'h14d == _T_54[9:0] ? px_buffer_333_r : _GEN_332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_334 = 10'h14e == _T_54[9:0] ? px_buffer_334_r : _GEN_333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_335 = 10'h14f == _T_54[9:0] ? px_buffer_335_r : _GEN_334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_336 = 10'h150 == _T_54[9:0] ? px_buffer_336_r : _GEN_335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_337 = 10'h151 == _T_54[9:0] ? px_buffer_337_r : _GEN_336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_338 = 10'h152 == _T_54[9:0] ? px_buffer_338_r : _GEN_337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_339 = 10'h153 == _T_54[9:0] ? px_buffer_339_r : _GEN_338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_340 = 10'h154 == _T_54[9:0] ? px_buffer_340_r : _GEN_339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_341 = 10'h155 == _T_54[9:0] ? px_buffer_341_r : _GEN_340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_342 = 10'h156 == _T_54[9:0] ? px_buffer_342_r : _GEN_341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_343 = 10'h157 == _T_54[9:0] ? px_buffer_343_r : _GEN_342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_344 = 10'h158 == _T_54[9:0] ? px_buffer_344_r : _GEN_343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_345 = 10'h159 == _T_54[9:0] ? px_buffer_345_r : _GEN_344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_346 = 10'h15a == _T_54[9:0] ? px_buffer_346_r : _GEN_345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_347 = 10'h15b == _T_54[9:0] ? px_buffer_347_r : _GEN_346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_348 = 10'h15c == _T_54[9:0] ? px_buffer_348_r : _GEN_347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_349 = 10'h15d == _T_54[9:0] ? px_buffer_349_r : _GEN_348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_350 = 10'h15e == _T_54[9:0] ? px_buffer_350_r : _GEN_349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_351 = 10'h15f == _T_54[9:0] ? px_buffer_351_r : _GEN_350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_352 = 10'h160 == _T_54[9:0] ? px_buffer_352_r : _GEN_351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_353 = 10'h161 == _T_54[9:0] ? px_buffer_353_r : _GEN_352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_354 = 10'h162 == _T_54[9:0] ? px_buffer_354_r : _GEN_353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_355 = 10'h163 == _T_54[9:0] ? px_buffer_355_r : _GEN_354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_356 = 10'h164 == _T_54[9:0] ? px_buffer_356_r : _GEN_355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_357 = 10'h165 == _T_54[9:0] ? px_buffer_357_r : _GEN_356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_358 = 10'h166 == _T_54[9:0] ? px_buffer_358_r : _GEN_357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_359 = 10'h167 == _T_54[9:0] ? px_buffer_359_r : _GEN_358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_360 = 10'h168 == _T_54[9:0] ? px_buffer_360_r : _GEN_359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_361 = 10'h169 == _T_54[9:0] ? px_buffer_361_r : _GEN_360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_362 = 10'h16a == _T_54[9:0] ? px_buffer_362_r : _GEN_361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_363 = 10'h16b == _T_54[9:0] ? px_buffer_363_r : _GEN_362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_364 = 10'h16c == _T_54[9:0] ? px_buffer_364_r : _GEN_363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_365 = 10'h16d == _T_54[9:0] ? px_buffer_365_r : _GEN_364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_366 = 10'h16e == _T_54[9:0] ? px_buffer_366_r : _GEN_365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_367 = 10'h16f == _T_54[9:0] ? px_buffer_367_r : _GEN_366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_368 = 10'h170 == _T_54[9:0] ? px_buffer_368_r : _GEN_367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_369 = 10'h171 == _T_54[9:0] ? px_buffer_369_r : _GEN_368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_370 = 10'h172 == _T_54[9:0] ? px_buffer_370_r : _GEN_369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_371 = 10'h173 == _T_54[9:0] ? px_buffer_371_r : _GEN_370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_372 = 10'h174 == _T_54[9:0] ? px_buffer_372_r : _GEN_371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_373 = 10'h175 == _T_54[9:0] ? px_buffer_373_r : _GEN_372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_374 = 10'h176 == _T_54[9:0] ? px_buffer_374_r : _GEN_373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_375 = 10'h177 == _T_54[9:0] ? px_buffer_375_r : _GEN_374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_376 = 10'h178 == _T_54[9:0] ? px_buffer_376_r : _GEN_375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_377 = 10'h179 == _T_54[9:0] ? px_buffer_377_r : _GEN_376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_378 = 10'h17a == _T_54[9:0] ? px_buffer_378_r : _GEN_377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_379 = 10'h17b == _T_54[9:0] ? px_buffer_379_r : _GEN_378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_380 = 10'h17c == _T_54[9:0] ? px_buffer_380_r : _GEN_379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_381 = 10'h17d == _T_54[9:0] ? px_buffer_381_r : _GEN_380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_382 = 10'h17e == _T_54[9:0] ? px_buffer_382_r : _GEN_381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_383 = 10'h17f == _T_54[9:0] ? px_buffer_383_r : _GEN_382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_384 = 10'h180 == _T_54[9:0] ? px_buffer_384_r : _GEN_383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_385 = 10'h181 == _T_54[9:0] ? px_buffer_385_r : _GEN_384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_386 = 10'h182 == _T_54[9:0] ? px_buffer_386_r : _GEN_385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_387 = 10'h183 == _T_54[9:0] ? px_buffer_387_r : _GEN_386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_388 = 10'h184 == _T_54[9:0] ? px_buffer_388_r : _GEN_387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_389 = 10'h185 == _T_54[9:0] ? px_buffer_389_r : _GEN_388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_390 = 10'h186 == _T_54[9:0] ? px_buffer_390_r : _GEN_389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_391 = 10'h187 == _T_54[9:0] ? px_buffer_391_r : _GEN_390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_392 = 10'h188 == _T_54[9:0] ? px_buffer_392_r : _GEN_391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_393 = 10'h189 == _T_54[9:0] ? px_buffer_393_r : _GEN_392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_394 = 10'h18a == _T_54[9:0] ? px_buffer_394_r : _GEN_393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_395 = 10'h18b == _T_54[9:0] ? px_buffer_395_r : _GEN_394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_396 = 10'h18c == _T_54[9:0] ? px_buffer_396_r : _GEN_395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_397 = 10'h18d == _T_54[9:0] ? px_buffer_397_r : _GEN_396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_398 = 10'h18e == _T_54[9:0] ? px_buffer_398_r : _GEN_397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_399 = 10'h18f == _T_54[9:0] ? px_buffer_399_r : _GEN_398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_400 = 10'h190 == _T_54[9:0] ? px_buffer_400_r : _GEN_399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_401 = 10'h191 == _T_54[9:0] ? px_buffer_401_r : _GEN_400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_402 = 10'h192 == _T_54[9:0] ? px_buffer_402_r : _GEN_401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_403 = 10'h193 == _T_54[9:0] ? px_buffer_403_r : _GEN_402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_404 = 10'h194 == _T_54[9:0] ? px_buffer_404_r : _GEN_403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_405 = 10'h195 == _T_54[9:0] ? px_buffer_405_r : _GEN_404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_406 = 10'h196 == _T_54[9:0] ? px_buffer_406_r : _GEN_405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_407 = 10'h197 == _T_54[9:0] ? px_buffer_407_r : _GEN_406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_408 = 10'h198 == _T_54[9:0] ? px_buffer_408_r : _GEN_407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_409 = 10'h199 == _T_54[9:0] ? px_buffer_409_r : _GEN_408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_410 = 10'h19a == _T_54[9:0] ? px_buffer_410_r : _GEN_409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_411 = 10'h19b == _T_54[9:0] ? px_buffer_411_r : _GEN_410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_412 = 10'h19c == _T_54[9:0] ? px_buffer_412_r : _GEN_411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_413 = 10'h19d == _T_54[9:0] ? px_buffer_413_r : _GEN_412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_414 = 10'h19e == _T_54[9:0] ? px_buffer_414_r : _GEN_413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_415 = 10'h19f == _T_54[9:0] ? px_buffer_415_r : _GEN_414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_416 = 10'h1a0 == _T_54[9:0] ? px_buffer_416_r : _GEN_415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_417 = 10'h1a1 == _T_54[9:0] ? px_buffer_417_r : _GEN_416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_418 = 10'h1a2 == _T_54[9:0] ? px_buffer_418_r : _GEN_417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_419 = 10'h1a3 == _T_54[9:0] ? px_buffer_419_r : _GEN_418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_420 = 10'h1a4 == _T_54[9:0] ? px_buffer_420_r : _GEN_419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_421 = 10'h1a5 == _T_54[9:0] ? px_buffer_421_r : _GEN_420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_422 = 10'h1a6 == _T_54[9:0] ? px_buffer_422_r : _GEN_421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_423 = 10'h1a7 == _T_54[9:0] ? px_buffer_423_r : _GEN_422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_424 = 10'h1a8 == _T_54[9:0] ? px_buffer_424_r : _GEN_423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_425 = 10'h1a9 == _T_54[9:0] ? px_buffer_425_r : _GEN_424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_426 = 10'h1aa == _T_54[9:0] ? px_buffer_426_r : _GEN_425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_427 = 10'h1ab == _T_54[9:0] ? px_buffer_427_r : _GEN_426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_428 = 10'h1ac == _T_54[9:0] ? px_buffer_428_r : _GEN_427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_429 = 10'h1ad == _T_54[9:0] ? px_buffer_429_r : _GEN_428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_430 = 10'h1ae == _T_54[9:0] ? px_buffer_430_r : _GEN_429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_431 = 10'h1af == _T_54[9:0] ? px_buffer_431_r : _GEN_430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_432 = 10'h1b0 == _T_54[9:0] ? px_buffer_432_r : _GEN_431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_433 = 10'h1b1 == _T_54[9:0] ? px_buffer_433_r : _GEN_432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_434 = 10'h1b2 == _T_54[9:0] ? px_buffer_434_r : _GEN_433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_435 = 10'h1b3 == _T_54[9:0] ? px_buffer_435_r : _GEN_434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_436 = 10'h1b4 == _T_54[9:0] ? px_buffer_436_r : _GEN_435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_437 = 10'h1b5 == _T_54[9:0] ? px_buffer_437_r : _GEN_436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_438 = 10'h1b6 == _T_54[9:0] ? px_buffer_438_r : _GEN_437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_439 = 10'h1b7 == _T_54[9:0] ? px_buffer_439_r : _GEN_438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_440 = 10'h1b8 == _T_54[9:0] ? px_buffer_440_r : _GEN_439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_441 = 10'h1b9 == _T_54[9:0] ? px_buffer_441_r : _GEN_440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_442 = 10'h1ba == _T_54[9:0] ? px_buffer_442_r : _GEN_441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_443 = 10'h1bb == _T_54[9:0] ? px_buffer_443_r : _GEN_442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_444 = 10'h1bc == _T_54[9:0] ? px_buffer_444_r : _GEN_443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_445 = 10'h1bd == _T_54[9:0] ? px_buffer_445_r : _GEN_444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_446 = 10'h1be == _T_54[9:0] ? px_buffer_446_r : _GEN_445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_447 = 10'h1bf == _T_54[9:0] ? px_buffer_447_r : _GEN_446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_448 = 10'h1c0 == _T_54[9:0] ? px_buffer_448_r : _GEN_447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_449 = 10'h1c1 == _T_54[9:0] ? px_buffer_449_r : _GEN_448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_450 = 10'h1c2 == _T_54[9:0] ? px_buffer_450_r : _GEN_449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_451 = 10'h1c3 == _T_54[9:0] ? px_buffer_451_r : _GEN_450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_452 = 10'h1c4 == _T_54[9:0] ? px_buffer_452_r : _GEN_451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_453 = 10'h1c5 == _T_54[9:0] ? px_buffer_453_r : _GEN_452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_454 = 10'h1c6 == _T_54[9:0] ? px_buffer_454_r : _GEN_453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_455 = 10'h1c7 == _T_54[9:0] ? px_buffer_455_r : _GEN_454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_456 = 10'h1c8 == _T_54[9:0] ? px_buffer_456_r : _GEN_455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_457 = 10'h1c9 == _T_54[9:0] ? px_buffer_457_r : _GEN_456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_458 = 10'h1ca == _T_54[9:0] ? px_buffer_458_r : _GEN_457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_459 = 10'h1cb == _T_54[9:0] ? px_buffer_459_r : _GEN_458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_460 = 10'h1cc == _T_54[9:0] ? px_buffer_460_r : _GEN_459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_461 = 10'h1cd == _T_54[9:0] ? px_buffer_461_r : _GEN_460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_462 = 10'h1ce == _T_54[9:0] ? px_buffer_462_r : _GEN_461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_463 = 10'h1cf == _T_54[9:0] ? px_buffer_463_r : _GEN_462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_464 = 10'h1d0 == _T_54[9:0] ? px_buffer_464_r : _GEN_463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_465 = 10'h1d1 == _T_54[9:0] ? px_buffer_465_r : _GEN_464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_466 = 10'h1d2 == _T_54[9:0] ? px_buffer_466_r : _GEN_465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_467 = 10'h1d3 == _T_54[9:0] ? px_buffer_467_r : _GEN_466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_468 = 10'h1d4 == _T_54[9:0] ? px_buffer_468_r : _GEN_467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_469 = 10'h1d5 == _T_54[9:0] ? px_buffer_469_r : _GEN_468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_470 = 10'h1d6 == _T_54[9:0] ? px_buffer_470_r : _GEN_469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_471 = 10'h1d7 == _T_54[9:0] ? px_buffer_471_r : _GEN_470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_472 = 10'h1d8 == _T_54[9:0] ? px_buffer_472_r : _GEN_471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_473 = 10'h1d9 == _T_54[9:0] ? px_buffer_473_r : _GEN_472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_474 = 10'h1da == _T_54[9:0] ? px_buffer_474_r : _GEN_473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_475 = 10'h1db == _T_54[9:0] ? px_buffer_475_r : _GEN_474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_476 = 10'h1dc == _T_54[9:0] ? px_buffer_476_r : _GEN_475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_477 = 10'h1dd == _T_54[9:0] ? px_buffer_477_r : _GEN_476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_478 = 10'h1de == _T_54[9:0] ? px_buffer_478_r : _GEN_477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_479 = 10'h1df == _T_54[9:0] ? px_buffer_479_r : _GEN_478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_480 = 10'h1e0 == _T_54[9:0] ? px_buffer_480_r : _GEN_479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_481 = 10'h1e1 == _T_54[9:0] ? px_buffer_481_r : _GEN_480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_482 = 10'h1e2 == _T_54[9:0] ? px_buffer_482_r : _GEN_481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_483 = 10'h1e3 == _T_54[9:0] ? px_buffer_483_r : _GEN_482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_484 = 10'h1e4 == _T_54[9:0] ? px_buffer_484_r : _GEN_483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_485 = 10'h1e5 == _T_54[9:0] ? px_buffer_485_r : _GEN_484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_486 = 10'h1e6 == _T_54[9:0] ? px_buffer_486_r : _GEN_485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_487 = 10'h1e7 == _T_54[9:0] ? px_buffer_487_r : _GEN_486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_488 = 10'h1e8 == _T_54[9:0] ? px_buffer_488_r : _GEN_487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_489 = 10'h1e9 == _T_54[9:0] ? px_buffer_489_r : _GEN_488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_490 = 10'h1ea == _T_54[9:0] ? px_buffer_490_r : _GEN_489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_491 = 10'h1eb == _T_54[9:0] ? px_buffer_491_r : _GEN_490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_492 = 10'h1ec == _T_54[9:0] ? px_buffer_492_r : _GEN_491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_493 = 10'h1ed == _T_54[9:0] ? px_buffer_493_r : _GEN_492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_494 = 10'h1ee == _T_54[9:0] ? px_buffer_494_r : _GEN_493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_495 = 10'h1ef == _T_54[9:0] ? px_buffer_495_r : _GEN_494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_496 = 10'h1f0 == _T_54[9:0] ? px_buffer_496_r : _GEN_495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_497 = 10'h1f1 == _T_54[9:0] ? px_buffer_497_r : _GEN_496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_498 = 10'h1f2 == _T_54[9:0] ? px_buffer_498_r : _GEN_497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_499 = 10'h1f3 == _T_54[9:0] ? px_buffer_499_r : _GEN_498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_500 = 10'h1f4 == _T_54[9:0] ? px_buffer_500_r : _GEN_499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_501 = 10'h1f5 == _T_54[9:0] ? px_buffer_501_r : _GEN_500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_502 = 10'h1f6 == _T_54[9:0] ? px_buffer_502_r : _GEN_501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_503 = 10'h1f7 == _T_54[9:0] ? px_buffer_503_r : _GEN_502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_504 = 10'h1f8 == _T_54[9:0] ? px_buffer_504_r : _GEN_503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_505 = 10'h1f9 == _T_54[9:0] ? px_buffer_505_r : _GEN_504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_506 = 10'h1fa == _T_54[9:0] ? px_buffer_506_r : _GEN_505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_507 = 10'h1fb == _T_54[9:0] ? px_buffer_507_r : _GEN_506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_508 = 10'h1fc == _T_54[9:0] ? px_buffer_508_r : _GEN_507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_509 = 10'h1fd == _T_54[9:0] ? px_buffer_509_r : _GEN_508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_510 = 10'h1fe == _T_54[9:0] ? px_buffer_510_r : _GEN_509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_511 = 10'h1ff == _T_54[9:0] ? px_buffer_511_r : _GEN_510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_512 = 10'h200 == _T_54[9:0] ? px_buffer_512_r : _GEN_511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_513 = 10'h201 == _T_54[9:0] ? px_buffer_513_r : _GEN_512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_514 = 10'h202 == _T_54[9:0] ? px_buffer_514_r : _GEN_513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_515 = 10'h203 == _T_54[9:0] ? px_buffer_515_r : _GEN_514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_516 = 10'h204 == _T_54[9:0] ? px_buffer_516_r : _GEN_515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_517 = 10'h205 == _T_54[9:0] ? px_buffer_517_r : _GEN_516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_518 = 10'h206 == _T_54[9:0] ? px_buffer_518_r : _GEN_517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_519 = 10'h207 == _T_54[9:0] ? px_buffer_519_r : _GEN_518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_520 = 10'h208 == _T_54[9:0] ? px_buffer_520_r : _GEN_519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_521 = 10'h209 == _T_54[9:0] ? px_buffer_521_r : _GEN_520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_522 = 10'h20a == _T_54[9:0] ? px_buffer_522_r : _GEN_521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_523 = 10'h20b == _T_54[9:0] ? px_buffer_523_r : _GEN_522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_524 = 10'h20c == _T_54[9:0] ? px_buffer_524_r : _GEN_523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_525 = 10'h20d == _T_54[9:0] ? px_buffer_525_r : _GEN_524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_526 = 10'h20e == _T_54[9:0] ? px_buffer_526_r : _GEN_525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_527 = 10'h20f == _T_54[9:0] ? px_buffer_527_r : _GEN_526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_528 = 10'h210 == _T_54[9:0] ? px_buffer_528_r : _GEN_527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_529 = 10'h211 == _T_54[9:0] ? px_buffer_529_r : _GEN_528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_530 = 10'h212 == _T_54[9:0] ? px_buffer_530_r : _GEN_529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_531 = 10'h213 == _T_54[9:0] ? px_buffer_531_r : _GEN_530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_532 = 10'h214 == _T_54[9:0] ? px_buffer_532_r : _GEN_531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_533 = 10'h215 == _T_54[9:0] ? px_buffer_533_r : _GEN_532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_534 = 10'h216 == _T_54[9:0] ? px_buffer_534_r : _GEN_533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_535 = 10'h217 == _T_54[9:0] ? px_buffer_535_r : _GEN_534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_536 = 10'h218 == _T_54[9:0] ? px_buffer_536_r : _GEN_535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_537 = 10'h219 == _T_54[9:0] ? px_buffer_537_r : _GEN_536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_538 = 10'h21a == _T_54[9:0] ? px_buffer_538_r : _GEN_537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_539 = 10'h21b == _T_54[9:0] ? px_buffer_539_r : _GEN_538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_540 = 10'h21c == _T_54[9:0] ? px_buffer_540_r : _GEN_539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_541 = 10'h21d == _T_54[9:0] ? px_buffer_541_r : _GEN_540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_542 = 10'h21e == _T_54[9:0] ? px_buffer_542_r : _GEN_541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_543 = 10'h21f == _T_54[9:0] ? px_buffer_543_r : _GEN_542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_544 = 10'h220 == _T_54[9:0] ? px_buffer_544_r : _GEN_543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_545 = 10'h221 == _T_54[9:0] ? px_buffer_545_r : _GEN_544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_546 = 10'h222 == _T_54[9:0] ? px_buffer_546_r : _GEN_545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_547 = 10'h223 == _T_54[9:0] ? px_buffer_547_r : _GEN_546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_548 = 10'h224 == _T_54[9:0] ? px_buffer_548_r : _GEN_547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_549 = 10'h225 == _T_54[9:0] ? px_buffer_549_r : _GEN_548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_550 = 10'h226 == _T_54[9:0] ? px_buffer_550_r : _GEN_549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_551 = 10'h227 == _T_54[9:0] ? px_buffer_551_r : _GEN_550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_552 = 10'h228 == _T_54[9:0] ? px_buffer_552_r : _GEN_551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_553 = 10'h229 == _T_54[9:0] ? px_buffer_553_r : _GEN_552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_554 = 10'h22a == _T_54[9:0] ? px_buffer_554_r : _GEN_553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_555 = 10'h22b == _T_54[9:0] ? px_buffer_555_r : _GEN_554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_556 = 10'h22c == _T_54[9:0] ? px_buffer_556_r : _GEN_555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_557 = 10'h22d == _T_54[9:0] ? px_buffer_557_r : _GEN_556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_558 = 10'h22e == _T_54[9:0] ? px_buffer_558_r : _GEN_557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_559 = 10'h22f == _T_54[9:0] ? px_buffer_559_r : _GEN_558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_560 = 10'h230 == _T_54[9:0] ? px_buffer_560_r : _GEN_559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_561 = 10'h231 == _T_54[9:0] ? px_buffer_561_r : _GEN_560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_562 = 10'h232 == _T_54[9:0] ? px_buffer_562_r : _GEN_561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_563 = 10'h233 == _T_54[9:0] ? px_buffer_563_r : _GEN_562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_564 = 10'h234 == _T_54[9:0] ? px_buffer_564_r : _GEN_563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_565 = 10'h235 == _T_54[9:0] ? px_buffer_565_r : _GEN_564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_566 = 10'h236 == _T_54[9:0] ? px_buffer_566_r : _GEN_565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_567 = 10'h237 == _T_54[9:0] ? px_buffer_567_r : _GEN_566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_568 = 10'h238 == _T_54[9:0] ? px_buffer_568_r : _GEN_567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_569 = 10'h239 == _T_54[9:0] ? px_buffer_569_r : _GEN_568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_570 = 10'h23a == _T_54[9:0] ? px_buffer_570_r : _GEN_569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_571 = 10'h23b == _T_54[9:0] ? px_buffer_571_r : _GEN_570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_572 = 10'h23c == _T_54[9:0] ? px_buffer_572_r : _GEN_571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_573 = 10'h23d == _T_54[9:0] ? px_buffer_573_r : _GEN_572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_574 = 10'h23e == _T_54[9:0] ? px_buffer_574_r : _GEN_573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_575 = 10'h23f == _T_54[9:0] ? px_buffer_575_r : _GEN_574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_576 = 10'h240 == _T_54[9:0] ? px_buffer_576_r : _GEN_575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_577 = 10'h241 == _T_54[9:0] ? px_buffer_577_r : _GEN_576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_578 = 10'h242 == _T_54[9:0] ? px_buffer_578_r : _GEN_577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_579 = 10'h243 == _T_54[9:0] ? px_buffer_579_r : _GEN_578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_580 = 10'h244 == _T_54[9:0] ? px_buffer_580_r : _GEN_579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_581 = 10'h245 == _T_54[9:0] ? px_buffer_581_r : _GEN_580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_582 = 10'h246 == _T_54[9:0] ? px_buffer_582_r : _GEN_581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_583 = 10'h247 == _T_54[9:0] ? px_buffer_583_r : _GEN_582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_584 = 10'h248 == _T_54[9:0] ? px_buffer_584_r : _GEN_583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_585 = 10'h249 == _T_54[9:0] ? px_buffer_585_r : _GEN_584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_586 = 10'h24a == _T_54[9:0] ? px_buffer_586_r : _GEN_585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_587 = 10'h24b == _T_54[9:0] ? px_buffer_587_r : _GEN_586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_588 = 10'h24c == _T_54[9:0] ? px_buffer_588_r : _GEN_587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_589 = 10'h24d == _T_54[9:0] ? px_buffer_589_r : _GEN_588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_590 = 10'h24e == _T_54[9:0] ? px_buffer_590_r : _GEN_589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_591 = 10'h24f == _T_54[9:0] ? px_buffer_591_r : _GEN_590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_592 = 10'h250 == _T_54[9:0] ? px_buffer_592_r : _GEN_591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_593 = 10'h251 == _T_54[9:0] ? px_buffer_593_r : _GEN_592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_594 = 10'h252 == _T_54[9:0] ? px_buffer_594_r : _GEN_593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_595 = 10'h253 == _T_54[9:0] ? px_buffer_595_r : _GEN_594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_596 = 10'h254 == _T_54[9:0] ? px_buffer_596_r : _GEN_595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_597 = 10'h255 == _T_54[9:0] ? px_buffer_597_r : _GEN_596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_598 = 10'h256 == _T_54[9:0] ? px_buffer_598_r : _GEN_597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_599 = 10'h257 == _T_54[9:0] ? px_buffer_599_r : _GEN_598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_600 = 10'h258 == _T_54[9:0] ? px_buffer_600_r : _GEN_599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_601 = 10'h259 == _T_54[9:0] ? px_buffer_601_r : _GEN_600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_602 = 10'h25a == _T_54[9:0] ? px_buffer_602_r : _GEN_601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_603 = 10'h25b == _T_54[9:0] ? px_buffer_603_r : _GEN_602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_604 = 10'h25c == _T_54[9:0] ? px_buffer_604_r : _GEN_603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_605 = 10'h25d == _T_54[9:0] ? px_buffer_605_r : _GEN_604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_606 = 10'h25e == _T_54[9:0] ? px_buffer_606_r : _GEN_605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_607 = 10'h25f == _T_54[9:0] ? px_buffer_607_r : _GEN_606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_608 = 10'h260 == _T_54[9:0] ? px_buffer_608_r : _GEN_607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_609 = 10'h261 == _T_54[9:0] ? px_buffer_609_r : _GEN_608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_610 = 10'h262 == _T_54[9:0] ? px_buffer_610_r : _GEN_609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_611 = 10'h263 == _T_54[9:0] ? px_buffer_611_r : _GEN_610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_612 = 10'h264 == _T_54[9:0] ? px_buffer_612_r : _GEN_611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_613 = 10'h265 == _T_54[9:0] ? px_buffer_613_r : _GEN_612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_614 = 10'h266 == _T_54[9:0] ? px_buffer_614_r : _GEN_613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_615 = 10'h267 == _T_54[9:0] ? px_buffer_615_r : _GEN_614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_616 = 10'h268 == _T_54[9:0] ? px_buffer_616_r : _GEN_615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_617 = 10'h269 == _T_54[9:0] ? px_buffer_617_r : _GEN_616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_618 = 10'h26a == _T_54[9:0] ? px_buffer_618_r : _GEN_617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_619 = 10'h26b == _T_54[9:0] ? px_buffer_619_r : _GEN_618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_620 = 10'h26c == _T_54[9:0] ? px_buffer_620_r : _GEN_619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_621 = 10'h26d == _T_54[9:0] ? px_buffer_621_r : _GEN_620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_622 = 10'h26e == _T_54[9:0] ? px_buffer_622_r : _GEN_621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_623 = 10'h26f == _T_54[9:0] ? px_buffer_623_r : _GEN_622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_624 = 10'h270 == _T_54[9:0] ? px_buffer_624_r : _GEN_623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_625 = 10'h271 == _T_54[9:0] ? px_buffer_625_r : _GEN_624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_626 = 10'h272 == _T_54[9:0] ? px_buffer_626_r : _GEN_625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_627 = 10'h273 == _T_54[9:0] ? px_buffer_627_r : _GEN_626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_628 = 10'h274 == _T_54[9:0] ? px_buffer_628_r : _GEN_627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_629 = 10'h275 == _T_54[9:0] ? px_buffer_629_r : _GEN_628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_630 = 10'h276 == _T_54[9:0] ? px_buffer_630_r : _GEN_629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_631 = 10'h277 == _T_54[9:0] ? px_buffer_631_r : _GEN_630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_632 = 10'h278 == _T_54[9:0] ? px_buffer_632_r : _GEN_631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_633 = 10'h279 == _T_54[9:0] ? px_buffer_633_r : _GEN_632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_634 = 10'h27a == _T_54[9:0] ? px_buffer_634_r : _GEN_633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_635 = 10'h27b == _T_54[9:0] ? px_buffer_635_r : _GEN_634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_636 = 10'h27c == _T_54[9:0] ? px_buffer_636_r : _GEN_635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_637 = 10'h27d == _T_54[9:0] ? px_buffer_637_r : _GEN_636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_638 = 10'h27e == _T_54[9:0] ? px_buffer_638_r : _GEN_637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_639 = 10'h27f == _T_54[9:0] ? px_buffer_639_r : _GEN_638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _T_57 = {1'h0,_GEN_639}; // @[EdgeDetect.scala 54:51]
  wire [8:0] _T_59 = {1'h0,io_px_in_r}; // @[EdgeDetect.scala 54:81]
  wire [8:0] _T_62 = $signed(_T_57) - $signed(_T_59); // @[EdgeDetect.scala 54:58]
  wire [7:0] _GEN_641 = 10'h1 == io_x[9:0] ? px_buffer_1_r : px_buffer_0_r; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_642 = 10'h2 == io_x[9:0] ? px_buffer_2_r : _GEN_641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_643 = 10'h3 == io_x[9:0] ? px_buffer_3_r : _GEN_642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_644 = 10'h4 == io_x[9:0] ? px_buffer_4_r : _GEN_643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_645 = 10'h5 == io_x[9:0] ? px_buffer_5_r : _GEN_644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_646 = 10'h6 == io_x[9:0] ? px_buffer_6_r : _GEN_645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_647 = 10'h7 == io_x[9:0] ? px_buffer_7_r : _GEN_646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_648 = 10'h8 == io_x[9:0] ? px_buffer_8_r : _GEN_647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_649 = 10'h9 == io_x[9:0] ? px_buffer_9_r : _GEN_648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_650 = 10'ha == io_x[9:0] ? px_buffer_10_r : _GEN_649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_651 = 10'hb == io_x[9:0] ? px_buffer_11_r : _GEN_650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_652 = 10'hc == io_x[9:0] ? px_buffer_12_r : _GEN_651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_653 = 10'hd == io_x[9:0] ? px_buffer_13_r : _GEN_652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_654 = 10'he == io_x[9:0] ? px_buffer_14_r : _GEN_653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_655 = 10'hf == io_x[9:0] ? px_buffer_15_r : _GEN_654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_656 = 10'h10 == io_x[9:0] ? px_buffer_16_r : _GEN_655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_657 = 10'h11 == io_x[9:0] ? px_buffer_17_r : _GEN_656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_658 = 10'h12 == io_x[9:0] ? px_buffer_18_r : _GEN_657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_659 = 10'h13 == io_x[9:0] ? px_buffer_19_r : _GEN_658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_660 = 10'h14 == io_x[9:0] ? px_buffer_20_r : _GEN_659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_661 = 10'h15 == io_x[9:0] ? px_buffer_21_r : _GEN_660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_662 = 10'h16 == io_x[9:0] ? px_buffer_22_r : _GEN_661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_663 = 10'h17 == io_x[9:0] ? px_buffer_23_r : _GEN_662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_664 = 10'h18 == io_x[9:0] ? px_buffer_24_r : _GEN_663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_665 = 10'h19 == io_x[9:0] ? px_buffer_25_r : _GEN_664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_666 = 10'h1a == io_x[9:0] ? px_buffer_26_r : _GEN_665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_667 = 10'h1b == io_x[9:0] ? px_buffer_27_r : _GEN_666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_668 = 10'h1c == io_x[9:0] ? px_buffer_28_r : _GEN_667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_669 = 10'h1d == io_x[9:0] ? px_buffer_29_r : _GEN_668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_670 = 10'h1e == io_x[9:0] ? px_buffer_30_r : _GEN_669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_671 = 10'h1f == io_x[9:0] ? px_buffer_31_r : _GEN_670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_672 = 10'h20 == io_x[9:0] ? px_buffer_32_r : _GEN_671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_673 = 10'h21 == io_x[9:0] ? px_buffer_33_r : _GEN_672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_674 = 10'h22 == io_x[9:0] ? px_buffer_34_r : _GEN_673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_675 = 10'h23 == io_x[9:0] ? px_buffer_35_r : _GEN_674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_676 = 10'h24 == io_x[9:0] ? px_buffer_36_r : _GEN_675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_677 = 10'h25 == io_x[9:0] ? px_buffer_37_r : _GEN_676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_678 = 10'h26 == io_x[9:0] ? px_buffer_38_r : _GEN_677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_679 = 10'h27 == io_x[9:0] ? px_buffer_39_r : _GEN_678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_680 = 10'h28 == io_x[9:0] ? px_buffer_40_r : _GEN_679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_681 = 10'h29 == io_x[9:0] ? px_buffer_41_r : _GEN_680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_682 = 10'h2a == io_x[9:0] ? px_buffer_42_r : _GEN_681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_683 = 10'h2b == io_x[9:0] ? px_buffer_43_r : _GEN_682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_684 = 10'h2c == io_x[9:0] ? px_buffer_44_r : _GEN_683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_685 = 10'h2d == io_x[9:0] ? px_buffer_45_r : _GEN_684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_686 = 10'h2e == io_x[9:0] ? px_buffer_46_r : _GEN_685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_687 = 10'h2f == io_x[9:0] ? px_buffer_47_r : _GEN_686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_688 = 10'h30 == io_x[9:0] ? px_buffer_48_r : _GEN_687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_689 = 10'h31 == io_x[9:0] ? px_buffer_49_r : _GEN_688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_690 = 10'h32 == io_x[9:0] ? px_buffer_50_r : _GEN_689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_691 = 10'h33 == io_x[9:0] ? px_buffer_51_r : _GEN_690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_692 = 10'h34 == io_x[9:0] ? px_buffer_52_r : _GEN_691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_693 = 10'h35 == io_x[9:0] ? px_buffer_53_r : _GEN_692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_694 = 10'h36 == io_x[9:0] ? px_buffer_54_r : _GEN_693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_695 = 10'h37 == io_x[9:0] ? px_buffer_55_r : _GEN_694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_696 = 10'h38 == io_x[9:0] ? px_buffer_56_r : _GEN_695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_697 = 10'h39 == io_x[9:0] ? px_buffer_57_r : _GEN_696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_698 = 10'h3a == io_x[9:0] ? px_buffer_58_r : _GEN_697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_699 = 10'h3b == io_x[9:0] ? px_buffer_59_r : _GEN_698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_700 = 10'h3c == io_x[9:0] ? px_buffer_60_r : _GEN_699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_701 = 10'h3d == io_x[9:0] ? px_buffer_61_r : _GEN_700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_702 = 10'h3e == io_x[9:0] ? px_buffer_62_r : _GEN_701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_703 = 10'h3f == io_x[9:0] ? px_buffer_63_r : _GEN_702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_704 = 10'h40 == io_x[9:0] ? px_buffer_64_r : _GEN_703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_705 = 10'h41 == io_x[9:0] ? px_buffer_65_r : _GEN_704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_706 = 10'h42 == io_x[9:0] ? px_buffer_66_r : _GEN_705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_707 = 10'h43 == io_x[9:0] ? px_buffer_67_r : _GEN_706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_708 = 10'h44 == io_x[9:0] ? px_buffer_68_r : _GEN_707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_709 = 10'h45 == io_x[9:0] ? px_buffer_69_r : _GEN_708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_710 = 10'h46 == io_x[9:0] ? px_buffer_70_r : _GEN_709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_711 = 10'h47 == io_x[9:0] ? px_buffer_71_r : _GEN_710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_712 = 10'h48 == io_x[9:0] ? px_buffer_72_r : _GEN_711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_713 = 10'h49 == io_x[9:0] ? px_buffer_73_r : _GEN_712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_714 = 10'h4a == io_x[9:0] ? px_buffer_74_r : _GEN_713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_715 = 10'h4b == io_x[9:0] ? px_buffer_75_r : _GEN_714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_716 = 10'h4c == io_x[9:0] ? px_buffer_76_r : _GEN_715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_717 = 10'h4d == io_x[9:0] ? px_buffer_77_r : _GEN_716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_718 = 10'h4e == io_x[9:0] ? px_buffer_78_r : _GEN_717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_719 = 10'h4f == io_x[9:0] ? px_buffer_79_r : _GEN_718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_720 = 10'h50 == io_x[9:0] ? px_buffer_80_r : _GEN_719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_721 = 10'h51 == io_x[9:0] ? px_buffer_81_r : _GEN_720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_722 = 10'h52 == io_x[9:0] ? px_buffer_82_r : _GEN_721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_723 = 10'h53 == io_x[9:0] ? px_buffer_83_r : _GEN_722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_724 = 10'h54 == io_x[9:0] ? px_buffer_84_r : _GEN_723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_725 = 10'h55 == io_x[9:0] ? px_buffer_85_r : _GEN_724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_726 = 10'h56 == io_x[9:0] ? px_buffer_86_r : _GEN_725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_727 = 10'h57 == io_x[9:0] ? px_buffer_87_r : _GEN_726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_728 = 10'h58 == io_x[9:0] ? px_buffer_88_r : _GEN_727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_729 = 10'h59 == io_x[9:0] ? px_buffer_89_r : _GEN_728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_730 = 10'h5a == io_x[9:0] ? px_buffer_90_r : _GEN_729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_731 = 10'h5b == io_x[9:0] ? px_buffer_91_r : _GEN_730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_732 = 10'h5c == io_x[9:0] ? px_buffer_92_r : _GEN_731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_733 = 10'h5d == io_x[9:0] ? px_buffer_93_r : _GEN_732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_734 = 10'h5e == io_x[9:0] ? px_buffer_94_r : _GEN_733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_735 = 10'h5f == io_x[9:0] ? px_buffer_95_r : _GEN_734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_736 = 10'h60 == io_x[9:0] ? px_buffer_96_r : _GEN_735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_737 = 10'h61 == io_x[9:0] ? px_buffer_97_r : _GEN_736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_738 = 10'h62 == io_x[9:0] ? px_buffer_98_r : _GEN_737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_739 = 10'h63 == io_x[9:0] ? px_buffer_99_r : _GEN_738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_740 = 10'h64 == io_x[9:0] ? px_buffer_100_r : _GEN_739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_741 = 10'h65 == io_x[9:0] ? px_buffer_101_r : _GEN_740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_742 = 10'h66 == io_x[9:0] ? px_buffer_102_r : _GEN_741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_743 = 10'h67 == io_x[9:0] ? px_buffer_103_r : _GEN_742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_744 = 10'h68 == io_x[9:0] ? px_buffer_104_r : _GEN_743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_745 = 10'h69 == io_x[9:0] ? px_buffer_105_r : _GEN_744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_746 = 10'h6a == io_x[9:0] ? px_buffer_106_r : _GEN_745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_747 = 10'h6b == io_x[9:0] ? px_buffer_107_r : _GEN_746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_748 = 10'h6c == io_x[9:0] ? px_buffer_108_r : _GEN_747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_749 = 10'h6d == io_x[9:0] ? px_buffer_109_r : _GEN_748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_750 = 10'h6e == io_x[9:0] ? px_buffer_110_r : _GEN_749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_751 = 10'h6f == io_x[9:0] ? px_buffer_111_r : _GEN_750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_752 = 10'h70 == io_x[9:0] ? px_buffer_112_r : _GEN_751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_753 = 10'h71 == io_x[9:0] ? px_buffer_113_r : _GEN_752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_754 = 10'h72 == io_x[9:0] ? px_buffer_114_r : _GEN_753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_755 = 10'h73 == io_x[9:0] ? px_buffer_115_r : _GEN_754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_756 = 10'h74 == io_x[9:0] ? px_buffer_116_r : _GEN_755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_757 = 10'h75 == io_x[9:0] ? px_buffer_117_r : _GEN_756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_758 = 10'h76 == io_x[9:0] ? px_buffer_118_r : _GEN_757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_759 = 10'h77 == io_x[9:0] ? px_buffer_119_r : _GEN_758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_760 = 10'h78 == io_x[9:0] ? px_buffer_120_r : _GEN_759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_761 = 10'h79 == io_x[9:0] ? px_buffer_121_r : _GEN_760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_762 = 10'h7a == io_x[9:0] ? px_buffer_122_r : _GEN_761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_763 = 10'h7b == io_x[9:0] ? px_buffer_123_r : _GEN_762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_764 = 10'h7c == io_x[9:0] ? px_buffer_124_r : _GEN_763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_765 = 10'h7d == io_x[9:0] ? px_buffer_125_r : _GEN_764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_766 = 10'h7e == io_x[9:0] ? px_buffer_126_r : _GEN_765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_767 = 10'h7f == io_x[9:0] ? px_buffer_127_r : _GEN_766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_768 = 10'h80 == io_x[9:0] ? px_buffer_128_r : _GEN_767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_769 = 10'h81 == io_x[9:0] ? px_buffer_129_r : _GEN_768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_770 = 10'h82 == io_x[9:0] ? px_buffer_130_r : _GEN_769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_771 = 10'h83 == io_x[9:0] ? px_buffer_131_r : _GEN_770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_772 = 10'h84 == io_x[9:0] ? px_buffer_132_r : _GEN_771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_773 = 10'h85 == io_x[9:0] ? px_buffer_133_r : _GEN_772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_774 = 10'h86 == io_x[9:0] ? px_buffer_134_r : _GEN_773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_775 = 10'h87 == io_x[9:0] ? px_buffer_135_r : _GEN_774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_776 = 10'h88 == io_x[9:0] ? px_buffer_136_r : _GEN_775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_777 = 10'h89 == io_x[9:0] ? px_buffer_137_r : _GEN_776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_778 = 10'h8a == io_x[9:0] ? px_buffer_138_r : _GEN_777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_779 = 10'h8b == io_x[9:0] ? px_buffer_139_r : _GEN_778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_780 = 10'h8c == io_x[9:0] ? px_buffer_140_r : _GEN_779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_781 = 10'h8d == io_x[9:0] ? px_buffer_141_r : _GEN_780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_782 = 10'h8e == io_x[9:0] ? px_buffer_142_r : _GEN_781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_783 = 10'h8f == io_x[9:0] ? px_buffer_143_r : _GEN_782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_784 = 10'h90 == io_x[9:0] ? px_buffer_144_r : _GEN_783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_785 = 10'h91 == io_x[9:0] ? px_buffer_145_r : _GEN_784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_786 = 10'h92 == io_x[9:0] ? px_buffer_146_r : _GEN_785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_787 = 10'h93 == io_x[9:0] ? px_buffer_147_r : _GEN_786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_788 = 10'h94 == io_x[9:0] ? px_buffer_148_r : _GEN_787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_789 = 10'h95 == io_x[9:0] ? px_buffer_149_r : _GEN_788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_790 = 10'h96 == io_x[9:0] ? px_buffer_150_r : _GEN_789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_791 = 10'h97 == io_x[9:0] ? px_buffer_151_r : _GEN_790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_792 = 10'h98 == io_x[9:0] ? px_buffer_152_r : _GEN_791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_793 = 10'h99 == io_x[9:0] ? px_buffer_153_r : _GEN_792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_794 = 10'h9a == io_x[9:0] ? px_buffer_154_r : _GEN_793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_795 = 10'h9b == io_x[9:0] ? px_buffer_155_r : _GEN_794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_796 = 10'h9c == io_x[9:0] ? px_buffer_156_r : _GEN_795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_797 = 10'h9d == io_x[9:0] ? px_buffer_157_r : _GEN_796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_798 = 10'h9e == io_x[9:0] ? px_buffer_158_r : _GEN_797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_799 = 10'h9f == io_x[9:0] ? px_buffer_159_r : _GEN_798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_800 = 10'ha0 == io_x[9:0] ? px_buffer_160_r : _GEN_799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_801 = 10'ha1 == io_x[9:0] ? px_buffer_161_r : _GEN_800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_802 = 10'ha2 == io_x[9:0] ? px_buffer_162_r : _GEN_801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_803 = 10'ha3 == io_x[9:0] ? px_buffer_163_r : _GEN_802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_804 = 10'ha4 == io_x[9:0] ? px_buffer_164_r : _GEN_803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_805 = 10'ha5 == io_x[9:0] ? px_buffer_165_r : _GEN_804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_806 = 10'ha6 == io_x[9:0] ? px_buffer_166_r : _GEN_805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_807 = 10'ha7 == io_x[9:0] ? px_buffer_167_r : _GEN_806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_808 = 10'ha8 == io_x[9:0] ? px_buffer_168_r : _GEN_807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_809 = 10'ha9 == io_x[9:0] ? px_buffer_169_r : _GEN_808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_810 = 10'haa == io_x[9:0] ? px_buffer_170_r : _GEN_809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_811 = 10'hab == io_x[9:0] ? px_buffer_171_r : _GEN_810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_812 = 10'hac == io_x[9:0] ? px_buffer_172_r : _GEN_811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_813 = 10'had == io_x[9:0] ? px_buffer_173_r : _GEN_812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_814 = 10'hae == io_x[9:0] ? px_buffer_174_r : _GEN_813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_815 = 10'haf == io_x[9:0] ? px_buffer_175_r : _GEN_814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_816 = 10'hb0 == io_x[9:0] ? px_buffer_176_r : _GEN_815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_817 = 10'hb1 == io_x[9:0] ? px_buffer_177_r : _GEN_816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_818 = 10'hb2 == io_x[9:0] ? px_buffer_178_r : _GEN_817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_819 = 10'hb3 == io_x[9:0] ? px_buffer_179_r : _GEN_818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_820 = 10'hb4 == io_x[9:0] ? px_buffer_180_r : _GEN_819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_821 = 10'hb5 == io_x[9:0] ? px_buffer_181_r : _GEN_820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_822 = 10'hb6 == io_x[9:0] ? px_buffer_182_r : _GEN_821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_823 = 10'hb7 == io_x[9:0] ? px_buffer_183_r : _GEN_822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_824 = 10'hb8 == io_x[9:0] ? px_buffer_184_r : _GEN_823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_825 = 10'hb9 == io_x[9:0] ? px_buffer_185_r : _GEN_824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_826 = 10'hba == io_x[9:0] ? px_buffer_186_r : _GEN_825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_827 = 10'hbb == io_x[9:0] ? px_buffer_187_r : _GEN_826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_828 = 10'hbc == io_x[9:0] ? px_buffer_188_r : _GEN_827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_829 = 10'hbd == io_x[9:0] ? px_buffer_189_r : _GEN_828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_830 = 10'hbe == io_x[9:0] ? px_buffer_190_r : _GEN_829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_831 = 10'hbf == io_x[9:0] ? px_buffer_191_r : _GEN_830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_832 = 10'hc0 == io_x[9:0] ? px_buffer_192_r : _GEN_831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_833 = 10'hc1 == io_x[9:0] ? px_buffer_193_r : _GEN_832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_834 = 10'hc2 == io_x[9:0] ? px_buffer_194_r : _GEN_833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_835 = 10'hc3 == io_x[9:0] ? px_buffer_195_r : _GEN_834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_836 = 10'hc4 == io_x[9:0] ? px_buffer_196_r : _GEN_835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_837 = 10'hc5 == io_x[9:0] ? px_buffer_197_r : _GEN_836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_838 = 10'hc6 == io_x[9:0] ? px_buffer_198_r : _GEN_837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_839 = 10'hc7 == io_x[9:0] ? px_buffer_199_r : _GEN_838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_840 = 10'hc8 == io_x[9:0] ? px_buffer_200_r : _GEN_839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_841 = 10'hc9 == io_x[9:0] ? px_buffer_201_r : _GEN_840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_842 = 10'hca == io_x[9:0] ? px_buffer_202_r : _GEN_841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_843 = 10'hcb == io_x[9:0] ? px_buffer_203_r : _GEN_842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_844 = 10'hcc == io_x[9:0] ? px_buffer_204_r : _GEN_843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_845 = 10'hcd == io_x[9:0] ? px_buffer_205_r : _GEN_844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_846 = 10'hce == io_x[9:0] ? px_buffer_206_r : _GEN_845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_847 = 10'hcf == io_x[9:0] ? px_buffer_207_r : _GEN_846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_848 = 10'hd0 == io_x[9:0] ? px_buffer_208_r : _GEN_847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_849 = 10'hd1 == io_x[9:0] ? px_buffer_209_r : _GEN_848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_850 = 10'hd2 == io_x[9:0] ? px_buffer_210_r : _GEN_849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_851 = 10'hd3 == io_x[9:0] ? px_buffer_211_r : _GEN_850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_852 = 10'hd4 == io_x[9:0] ? px_buffer_212_r : _GEN_851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_853 = 10'hd5 == io_x[9:0] ? px_buffer_213_r : _GEN_852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_854 = 10'hd6 == io_x[9:0] ? px_buffer_214_r : _GEN_853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_855 = 10'hd7 == io_x[9:0] ? px_buffer_215_r : _GEN_854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_856 = 10'hd8 == io_x[9:0] ? px_buffer_216_r : _GEN_855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_857 = 10'hd9 == io_x[9:0] ? px_buffer_217_r : _GEN_856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_858 = 10'hda == io_x[9:0] ? px_buffer_218_r : _GEN_857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_859 = 10'hdb == io_x[9:0] ? px_buffer_219_r : _GEN_858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_860 = 10'hdc == io_x[9:0] ? px_buffer_220_r : _GEN_859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_861 = 10'hdd == io_x[9:0] ? px_buffer_221_r : _GEN_860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_862 = 10'hde == io_x[9:0] ? px_buffer_222_r : _GEN_861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_863 = 10'hdf == io_x[9:0] ? px_buffer_223_r : _GEN_862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_864 = 10'he0 == io_x[9:0] ? px_buffer_224_r : _GEN_863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_865 = 10'he1 == io_x[9:0] ? px_buffer_225_r : _GEN_864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_866 = 10'he2 == io_x[9:0] ? px_buffer_226_r : _GEN_865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_867 = 10'he3 == io_x[9:0] ? px_buffer_227_r : _GEN_866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_868 = 10'he4 == io_x[9:0] ? px_buffer_228_r : _GEN_867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_869 = 10'he5 == io_x[9:0] ? px_buffer_229_r : _GEN_868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_870 = 10'he6 == io_x[9:0] ? px_buffer_230_r : _GEN_869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_871 = 10'he7 == io_x[9:0] ? px_buffer_231_r : _GEN_870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_872 = 10'he8 == io_x[9:0] ? px_buffer_232_r : _GEN_871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_873 = 10'he9 == io_x[9:0] ? px_buffer_233_r : _GEN_872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_874 = 10'hea == io_x[9:0] ? px_buffer_234_r : _GEN_873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_875 = 10'heb == io_x[9:0] ? px_buffer_235_r : _GEN_874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_876 = 10'hec == io_x[9:0] ? px_buffer_236_r : _GEN_875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_877 = 10'hed == io_x[9:0] ? px_buffer_237_r : _GEN_876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_878 = 10'hee == io_x[9:0] ? px_buffer_238_r : _GEN_877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_879 = 10'hef == io_x[9:0] ? px_buffer_239_r : _GEN_878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_880 = 10'hf0 == io_x[9:0] ? px_buffer_240_r : _GEN_879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_881 = 10'hf1 == io_x[9:0] ? px_buffer_241_r : _GEN_880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_882 = 10'hf2 == io_x[9:0] ? px_buffer_242_r : _GEN_881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_883 = 10'hf3 == io_x[9:0] ? px_buffer_243_r : _GEN_882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_884 = 10'hf4 == io_x[9:0] ? px_buffer_244_r : _GEN_883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_885 = 10'hf5 == io_x[9:0] ? px_buffer_245_r : _GEN_884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_886 = 10'hf6 == io_x[9:0] ? px_buffer_246_r : _GEN_885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_887 = 10'hf7 == io_x[9:0] ? px_buffer_247_r : _GEN_886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_888 = 10'hf8 == io_x[9:0] ? px_buffer_248_r : _GEN_887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_889 = 10'hf9 == io_x[9:0] ? px_buffer_249_r : _GEN_888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_890 = 10'hfa == io_x[9:0] ? px_buffer_250_r : _GEN_889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_891 = 10'hfb == io_x[9:0] ? px_buffer_251_r : _GEN_890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_892 = 10'hfc == io_x[9:0] ? px_buffer_252_r : _GEN_891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_893 = 10'hfd == io_x[9:0] ? px_buffer_253_r : _GEN_892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_894 = 10'hfe == io_x[9:0] ? px_buffer_254_r : _GEN_893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_895 = 10'hff == io_x[9:0] ? px_buffer_255_r : _GEN_894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_896 = 10'h100 == io_x[9:0] ? px_buffer_256_r : _GEN_895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_897 = 10'h101 == io_x[9:0] ? px_buffer_257_r : _GEN_896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_898 = 10'h102 == io_x[9:0] ? px_buffer_258_r : _GEN_897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_899 = 10'h103 == io_x[9:0] ? px_buffer_259_r : _GEN_898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_900 = 10'h104 == io_x[9:0] ? px_buffer_260_r : _GEN_899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_901 = 10'h105 == io_x[9:0] ? px_buffer_261_r : _GEN_900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_902 = 10'h106 == io_x[9:0] ? px_buffer_262_r : _GEN_901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_903 = 10'h107 == io_x[9:0] ? px_buffer_263_r : _GEN_902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_904 = 10'h108 == io_x[9:0] ? px_buffer_264_r : _GEN_903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_905 = 10'h109 == io_x[9:0] ? px_buffer_265_r : _GEN_904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_906 = 10'h10a == io_x[9:0] ? px_buffer_266_r : _GEN_905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_907 = 10'h10b == io_x[9:0] ? px_buffer_267_r : _GEN_906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_908 = 10'h10c == io_x[9:0] ? px_buffer_268_r : _GEN_907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_909 = 10'h10d == io_x[9:0] ? px_buffer_269_r : _GEN_908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_910 = 10'h10e == io_x[9:0] ? px_buffer_270_r : _GEN_909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_911 = 10'h10f == io_x[9:0] ? px_buffer_271_r : _GEN_910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_912 = 10'h110 == io_x[9:0] ? px_buffer_272_r : _GEN_911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_913 = 10'h111 == io_x[9:0] ? px_buffer_273_r : _GEN_912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_914 = 10'h112 == io_x[9:0] ? px_buffer_274_r : _GEN_913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_915 = 10'h113 == io_x[9:0] ? px_buffer_275_r : _GEN_914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_916 = 10'h114 == io_x[9:0] ? px_buffer_276_r : _GEN_915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_917 = 10'h115 == io_x[9:0] ? px_buffer_277_r : _GEN_916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_918 = 10'h116 == io_x[9:0] ? px_buffer_278_r : _GEN_917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_919 = 10'h117 == io_x[9:0] ? px_buffer_279_r : _GEN_918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_920 = 10'h118 == io_x[9:0] ? px_buffer_280_r : _GEN_919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_921 = 10'h119 == io_x[9:0] ? px_buffer_281_r : _GEN_920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_922 = 10'h11a == io_x[9:0] ? px_buffer_282_r : _GEN_921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_923 = 10'h11b == io_x[9:0] ? px_buffer_283_r : _GEN_922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_924 = 10'h11c == io_x[9:0] ? px_buffer_284_r : _GEN_923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_925 = 10'h11d == io_x[9:0] ? px_buffer_285_r : _GEN_924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_926 = 10'h11e == io_x[9:0] ? px_buffer_286_r : _GEN_925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_927 = 10'h11f == io_x[9:0] ? px_buffer_287_r : _GEN_926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_928 = 10'h120 == io_x[9:0] ? px_buffer_288_r : _GEN_927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_929 = 10'h121 == io_x[9:0] ? px_buffer_289_r : _GEN_928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_930 = 10'h122 == io_x[9:0] ? px_buffer_290_r : _GEN_929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_931 = 10'h123 == io_x[9:0] ? px_buffer_291_r : _GEN_930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_932 = 10'h124 == io_x[9:0] ? px_buffer_292_r : _GEN_931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_933 = 10'h125 == io_x[9:0] ? px_buffer_293_r : _GEN_932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_934 = 10'h126 == io_x[9:0] ? px_buffer_294_r : _GEN_933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_935 = 10'h127 == io_x[9:0] ? px_buffer_295_r : _GEN_934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_936 = 10'h128 == io_x[9:0] ? px_buffer_296_r : _GEN_935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_937 = 10'h129 == io_x[9:0] ? px_buffer_297_r : _GEN_936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_938 = 10'h12a == io_x[9:0] ? px_buffer_298_r : _GEN_937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_939 = 10'h12b == io_x[9:0] ? px_buffer_299_r : _GEN_938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_940 = 10'h12c == io_x[9:0] ? px_buffer_300_r : _GEN_939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_941 = 10'h12d == io_x[9:0] ? px_buffer_301_r : _GEN_940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_942 = 10'h12e == io_x[9:0] ? px_buffer_302_r : _GEN_941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_943 = 10'h12f == io_x[9:0] ? px_buffer_303_r : _GEN_942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_944 = 10'h130 == io_x[9:0] ? px_buffer_304_r : _GEN_943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_945 = 10'h131 == io_x[9:0] ? px_buffer_305_r : _GEN_944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_946 = 10'h132 == io_x[9:0] ? px_buffer_306_r : _GEN_945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_947 = 10'h133 == io_x[9:0] ? px_buffer_307_r : _GEN_946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_948 = 10'h134 == io_x[9:0] ? px_buffer_308_r : _GEN_947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_949 = 10'h135 == io_x[9:0] ? px_buffer_309_r : _GEN_948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_950 = 10'h136 == io_x[9:0] ? px_buffer_310_r : _GEN_949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_951 = 10'h137 == io_x[9:0] ? px_buffer_311_r : _GEN_950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_952 = 10'h138 == io_x[9:0] ? px_buffer_312_r : _GEN_951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_953 = 10'h139 == io_x[9:0] ? px_buffer_313_r : _GEN_952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_954 = 10'h13a == io_x[9:0] ? px_buffer_314_r : _GEN_953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_955 = 10'h13b == io_x[9:0] ? px_buffer_315_r : _GEN_954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_956 = 10'h13c == io_x[9:0] ? px_buffer_316_r : _GEN_955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_957 = 10'h13d == io_x[9:0] ? px_buffer_317_r : _GEN_956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_958 = 10'h13e == io_x[9:0] ? px_buffer_318_r : _GEN_957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_959 = 10'h13f == io_x[9:0] ? px_buffer_319_r : _GEN_958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_960 = 10'h140 == io_x[9:0] ? px_buffer_320_r : _GEN_959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_961 = 10'h141 == io_x[9:0] ? px_buffer_321_r : _GEN_960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_962 = 10'h142 == io_x[9:0] ? px_buffer_322_r : _GEN_961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_963 = 10'h143 == io_x[9:0] ? px_buffer_323_r : _GEN_962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_964 = 10'h144 == io_x[9:0] ? px_buffer_324_r : _GEN_963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_965 = 10'h145 == io_x[9:0] ? px_buffer_325_r : _GEN_964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_966 = 10'h146 == io_x[9:0] ? px_buffer_326_r : _GEN_965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_967 = 10'h147 == io_x[9:0] ? px_buffer_327_r : _GEN_966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_968 = 10'h148 == io_x[9:0] ? px_buffer_328_r : _GEN_967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_969 = 10'h149 == io_x[9:0] ? px_buffer_329_r : _GEN_968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_970 = 10'h14a == io_x[9:0] ? px_buffer_330_r : _GEN_969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_971 = 10'h14b == io_x[9:0] ? px_buffer_331_r : _GEN_970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_972 = 10'h14c == io_x[9:0] ? px_buffer_332_r : _GEN_971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_973 = 10'h14d == io_x[9:0] ? px_buffer_333_r : _GEN_972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_974 = 10'h14e == io_x[9:0] ? px_buffer_334_r : _GEN_973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_975 = 10'h14f == io_x[9:0] ? px_buffer_335_r : _GEN_974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_976 = 10'h150 == io_x[9:0] ? px_buffer_336_r : _GEN_975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_977 = 10'h151 == io_x[9:0] ? px_buffer_337_r : _GEN_976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_978 = 10'h152 == io_x[9:0] ? px_buffer_338_r : _GEN_977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_979 = 10'h153 == io_x[9:0] ? px_buffer_339_r : _GEN_978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_980 = 10'h154 == io_x[9:0] ? px_buffer_340_r : _GEN_979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_981 = 10'h155 == io_x[9:0] ? px_buffer_341_r : _GEN_980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_982 = 10'h156 == io_x[9:0] ? px_buffer_342_r : _GEN_981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_983 = 10'h157 == io_x[9:0] ? px_buffer_343_r : _GEN_982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_984 = 10'h158 == io_x[9:0] ? px_buffer_344_r : _GEN_983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_985 = 10'h159 == io_x[9:0] ? px_buffer_345_r : _GEN_984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_986 = 10'h15a == io_x[9:0] ? px_buffer_346_r : _GEN_985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_987 = 10'h15b == io_x[9:0] ? px_buffer_347_r : _GEN_986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_988 = 10'h15c == io_x[9:0] ? px_buffer_348_r : _GEN_987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_989 = 10'h15d == io_x[9:0] ? px_buffer_349_r : _GEN_988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_990 = 10'h15e == io_x[9:0] ? px_buffer_350_r : _GEN_989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_991 = 10'h15f == io_x[9:0] ? px_buffer_351_r : _GEN_990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_992 = 10'h160 == io_x[9:0] ? px_buffer_352_r : _GEN_991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_993 = 10'h161 == io_x[9:0] ? px_buffer_353_r : _GEN_992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_994 = 10'h162 == io_x[9:0] ? px_buffer_354_r : _GEN_993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_995 = 10'h163 == io_x[9:0] ? px_buffer_355_r : _GEN_994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_996 = 10'h164 == io_x[9:0] ? px_buffer_356_r : _GEN_995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_997 = 10'h165 == io_x[9:0] ? px_buffer_357_r : _GEN_996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_998 = 10'h166 == io_x[9:0] ? px_buffer_358_r : _GEN_997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_999 = 10'h167 == io_x[9:0] ? px_buffer_359_r : _GEN_998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1000 = 10'h168 == io_x[9:0] ? px_buffer_360_r : _GEN_999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1001 = 10'h169 == io_x[9:0] ? px_buffer_361_r : _GEN_1000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1002 = 10'h16a == io_x[9:0] ? px_buffer_362_r : _GEN_1001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1003 = 10'h16b == io_x[9:0] ? px_buffer_363_r : _GEN_1002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1004 = 10'h16c == io_x[9:0] ? px_buffer_364_r : _GEN_1003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1005 = 10'h16d == io_x[9:0] ? px_buffer_365_r : _GEN_1004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1006 = 10'h16e == io_x[9:0] ? px_buffer_366_r : _GEN_1005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1007 = 10'h16f == io_x[9:0] ? px_buffer_367_r : _GEN_1006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1008 = 10'h170 == io_x[9:0] ? px_buffer_368_r : _GEN_1007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1009 = 10'h171 == io_x[9:0] ? px_buffer_369_r : _GEN_1008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1010 = 10'h172 == io_x[9:0] ? px_buffer_370_r : _GEN_1009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1011 = 10'h173 == io_x[9:0] ? px_buffer_371_r : _GEN_1010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1012 = 10'h174 == io_x[9:0] ? px_buffer_372_r : _GEN_1011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1013 = 10'h175 == io_x[9:0] ? px_buffer_373_r : _GEN_1012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1014 = 10'h176 == io_x[9:0] ? px_buffer_374_r : _GEN_1013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1015 = 10'h177 == io_x[9:0] ? px_buffer_375_r : _GEN_1014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1016 = 10'h178 == io_x[9:0] ? px_buffer_376_r : _GEN_1015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1017 = 10'h179 == io_x[9:0] ? px_buffer_377_r : _GEN_1016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1018 = 10'h17a == io_x[9:0] ? px_buffer_378_r : _GEN_1017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1019 = 10'h17b == io_x[9:0] ? px_buffer_379_r : _GEN_1018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1020 = 10'h17c == io_x[9:0] ? px_buffer_380_r : _GEN_1019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1021 = 10'h17d == io_x[9:0] ? px_buffer_381_r : _GEN_1020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1022 = 10'h17e == io_x[9:0] ? px_buffer_382_r : _GEN_1021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1023 = 10'h17f == io_x[9:0] ? px_buffer_383_r : _GEN_1022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1024 = 10'h180 == io_x[9:0] ? px_buffer_384_r : _GEN_1023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1025 = 10'h181 == io_x[9:0] ? px_buffer_385_r : _GEN_1024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1026 = 10'h182 == io_x[9:0] ? px_buffer_386_r : _GEN_1025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1027 = 10'h183 == io_x[9:0] ? px_buffer_387_r : _GEN_1026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1028 = 10'h184 == io_x[9:0] ? px_buffer_388_r : _GEN_1027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1029 = 10'h185 == io_x[9:0] ? px_buffer_389_r : _GEN_1028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1030 = 10'h186 == io_x[9:0] ? px_buffer_390_r : _GEN_1029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1031 = 10'h187 == io_x[9:0] ? px_buffer_391_r : _GEN_1030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1032 = 10'h188 == io_x[9:0] ? px_buffer_392_r : _GEN_1031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1033 = 10'h189 == io_x[9:0] ? px_buffer_393_r : _GEN_1032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1034 = 10'h18a == io_x[9:0] ? px_buffer_394_r : _GEN_1033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1035 = 10'h18b == io_x[9:0] ? px_buffer_395_r : _GEN_1034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1036 = 10'h18c == io_x[9:0] ? px_buffer_396_r : _GEN_1035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1037 = 10'h18d == io_x[9:0] ? px_buffer_397_r : _GEN_1036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1038 = 10'h18e == io_x[9:0] ? px_buffer_398_r : _GEN_1037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1039 = 10'h18f == io_x[9:0] ? px_buffer_399_r : _GEN_1038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1040 = 10'h190 == io_x[9:0] ? px_buffer_400_r : _GEN_1039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1041 = 10'h191 == io_x[9:0] ? px_buffer_401_r : _GEN_1040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1042 = 10'h192 == io_x[9:0] ? px_buffer_402_r : _GEN_1041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1043 = 10'h193 == io_x[9:0] ? px_buffer_403_r : _GEN_1042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1044 = 10'h194 == io_x[9:0] ? px_buffer_404_r : _GEN_1043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1045 = 10'h195 == io_x[9:0] ? px_buffer_405_r : _GEN_1044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1046 = 10'h196 == io_x[9:0] ? px_buffer_406_r : _GEN_1045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1047 = 10'h197 == io_x[9:0] ? px_buffer_407_r : _GEN_1046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1048 = 10'h198 == io_x[9:0] ? px_buffer_408_r : _GEN_1047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1049 = 10'h199 == io_x[9:0] ? px_buffer_409_r : _GEN_1048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1050 = 10'h19a == io_x[9:0] ? px_buffer_410_r : _GEN_1049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1051 = 10'h19b == io_x[9:0] ? px_buffer_411_r : _GEN_1050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1052 = 10'h19c == io_x[9:0] ? px_buffer_412_r : _GEN_1051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1053 = 10'h19d == io_x[9:0] ? px_buffer_413_r : _GEN_1052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1054 = 10'h19e == io_x[9:0] ? px_buffer_414_r : _GEN_1053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1055 = 10'h19f == io_x[9:0] ? px_buffer_415_r : _GEN_1054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1056 = 10'h1a0 == io_x[9:0] ? px_buffer_416_r : _GEN_1055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1057 = 10'h1a1 == io_x[9:0] ? px_buffer_417_r : _GEN_1056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1058 = 10'h1a2 == io_x[9:0] ? px_buffer_418_r : _GEN_1057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1059 = 10'h1a3 == io_x[9:0] ? px_buffer_419_r : _GEN_1058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1060 = 10'h1a4 == io_x[9:0] ? px_buffer_420_r : _GEN_1059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1061 = 10'h1a5 == io_x[9:0] ? px_buffer_421_r : _GEN_1060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1062 = 10'h1a6 == io_x[9:0] ? px_buffer_422_r : _GEN_1061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1063 = 10'h1a7 == io_x[9:0] ? px_buffer_423_r : _GEN_1062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1064 = 10'h1a8 == io_x[9:0] ? px_buffer_424_r : _GEN_1063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1065 = 10'h1a9 == io_x[9:0] ? px_buffer_425_r : _GEN_1064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1066 = 10'h1aa == io_x[9:0] ? px_buffer_426_r : _GEN_1065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1067 = 10'h1ab == io_x[9:0] ? px_buffer_427_r : _GEN_1066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1068 = 10'h1ac == io_x[9:0] ? px_buffer_428_r : _GEN_1067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1069 = 10'h1ad == io_x[9:0] ? px_buffer_429_r : _GEN_1068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1070 = 10'h1ae == io_x[9:0] ? px_buffer_430_r : _GEN_1069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1071 = 10'h1af == io_x[9:0] ? px_buffer_431_r : _GEN_1070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1072 = 10'h1b0 == io_x[9:0] ? px_buffer_432_r : _GEN_1071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1073 = 10'h1b1 == io_x[9:0] ? px_buffer_433_r : _GEN_1072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1074 = 10'h1b2 == io_x[9:0] ? px_buffer_434_r : _GEN_1073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1075 = 10'h1b3 == io_x[9:0] ? px_buffer_435_r : _GEN_1074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1076 = 10'h1b4 == io_x[9:0] ? px_buffer_436_r : _GEN_1075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1077 = 10'h1b5 == io_x[9:0] ? px_buffer_437_r : _GEN_1076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1078 = 10'h1b6 == io_x[9:0] ? px_buffer_438_r : _GEN_1077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1079 = 10'h1b7 == io_x[9:0] ? px_buffer_439_r : _GEN_1078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1080 = 10'h1b8 == io_x[9:0] ? px_buffer_440_r : _GEN_1079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1081 = 10'h1b9 == io_x[9:0] ? px_buffer_441_r : _GEN_1080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1082 = 10'h1ba == io_x[9:0] ? px_buffer_442_r : _GEN_1081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1083 = 10'h1bb == io_x[9:0] ? px_buffer_443_r : _GEN_1082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1084 = 10'h1bc == io_x[9:0] ? px_buffer_444_r : _GEN_1083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1085 = 10'h1bd == io_x[9:0] ? px_buffer_445_r : _GEN_1084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1086 = 10'h1be == io_x[9:0] ? px_buffer_446_r : _GEN_1085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1087 = 10'h1bf == io_x[9:0] ? px_buffer_447_r : _GEN_1086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1088 = 10'h1c0 == io_x[9:0] ? px_buffer_448_r : _GEN_1087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1089 = 10'h1c1 == io_x[9:0] ? px_buffer_449_r : _GEN_1088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1090 = 10'h1c2 == io_x[9:0] ? px_buffer_450_r : _GEN_1089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1091 = 10'h1c3 == io_x[9:0] ? px_buffer_451_r : _GEN_1090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1092 = 10'h1c4 == io_x[9:0] ? px_buffer_452_r : _GEN_1091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1093 = 10'h1c5 == io_x[9:0] ? px_buffer_453_r : _GEN_1092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1094 = 10'h1c6 == io_x[9:0] ? px_buffer_454_r : _GEN_1093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1095 = 10'h1c7 == io_x[9:0] ? px_buffer_455_r : _GEN_1094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1096 = 10'h1c8 == io_x[9:0] ? px_buffer_456_r : _GEN_1095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1097 = 10'h1c9 == io_x[9:0] ? px_buffer_457_r : _GEN_1096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1098 = 10'h1ca == io_x[9:0] ? px_buffer_458_r : _GEN_1097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1099 = 10'h1cb == io_x[9:0] ? px_buffer_459_r : _GEN_1098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1100 = 10'h1cc == io_x[9:0] ? px_buffer_460_r : _GEN_1099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1101 = 10'h1cd == io_x[9:0] ? px_buffer_461_r : _GEN_1100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1102 = 10'h1ce == io_x[9:0] ? px_buffer_462_r : _GEN_1101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1103 = 10'h1cf == io_x[9:0] ? px_buffer_463_r : _GEN_1102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1104 = 10'h1d0 == io_x[9:0] ? px_buffer_464_r : _GEN_1103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1105 = 10'h1d1 == io_x[9:0] ? px_buffer_465_r : _GEN_1104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1106 = 10'h1d2 == io_x[9:0] ? px_buffer_466_r : _GEN_1105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1107 = 10'h1d3 == io_x[9:0] ? px_buffer_467_r : _GEN_1106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1108 = 10'h1d4 == io_x[9:0] ? px_buffer_468_r : _GEN_1107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1109 = 10'h1d5 == io_x[9:0] ? px_buffer_469_r : _GEN_1108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1110 = 10'h1d6 == io_x[9:0] ? px_buffer_470_r : _GEN_1109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1111 = 10'h1d7 == io_x[9:0] ? px_buffer_471_r : _GEN_1110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1112 = 10'h1d8 == io_x[9:0] ? px_buffer_472_r : _GEN_1111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1113 = 10'h1d9 == io_x[9:0] ? px_buffer_473_r : _GEN_1112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1114 = 10'h1da == io_x[9:0] ? px_buffer_474_r : _GEN_1113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1115 = 10'h1db == io_x[9:0] ? px_buffer_475_r : _GEN_1114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1116 = 10'h1dc == io_x[9:0] ? px_buffer_476_r : _GEN_1115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1117 = 10'h1dd == io_x[9:0] ? px_buffer_477_r : _GEN_1116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1118 = 10'h1de == io_x[9:0] ? px_buffer_478_r : _GEN_1117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1119 = 10'h1df == io_x[9:0] ? px_buffer_479_r : _GEN_1118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1120 = 10'h1e0 == io_x[9:0] ? px_buffer_480_r : _GEN_1119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1121 = 10'h1e1 == io_x[9:0] ? px_buffer_481_r : _GEN_1120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1122 = 10'h1e2 == io_x[9:0] ? px_buffer_482_r : _GEN_1121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1123 = 10'h1e3 == io_x[9:0] ? px_buffer_483_r : _GEN_1122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1124 = 10'h1e4 == io_x[9:0] ? px_buffer_484_r : _GEN_1123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1125 = 10'h1e5 == io_x[9:0] ? px_buffer_485_r : _GEN_1124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1126 = 10'h1e6 == io_x[9:0] ? px_buffer_486_r : _GEN_1125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1127 = 10'h1e7 == io_x[9:0] ? px_buffer_487_r : _GEN_1126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1128 = 10'h1e8 == io_x[9:0] ? px_buffer_488_r : _GEN_1127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1129 = 10'h1e9 == io_x[9:0] ? px_buffer_489_r : _GEN_1128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1130 = 10'h1ea == io_x[9:0] ? px_buffer_490_r : _GEN_1129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1131 = 10'h1eb == io_x[9:0] ? px_buffer_491_r : _GEN_1130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1132 = 10'h1ec == io_x[9:0] ? px_buffer_492_r : _GEN_1131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1133 = 10'h1ed == io_x[9:0] ? px_buffer_493_r : _GEN_1132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1134 = 10'h1ee == io_x[9:0] ? px_buffer_494_r : _GEN_1133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1135 = 10'h1ef == io_x[9:0] ? px_buffer_495_r : _GEN_1134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1136 = 10'h1f0 == io_x[9:0] ? px_buffer_496_r : _GEN_1135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1137 = 10'h1f1 == io_x[9:0] ? px_buffer_497_r : _GEN_1136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1138 = 10'h1f2 == io_x[9:0] ? px_buffer_498_r : _GEN_1137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1139 = 10'h1f3 == io_x[9:0] ? px_buffer_499_r : _GEN_1138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1140 = 10'h1f4 == io_x[9:0] ? px_buffer_500_r : _GEN_1139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1141 = 10'h1f5 == io_x[9:0] ? px_buffer_501_r : _GEN_1140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1142 = 10'h1f6 == io_x[9:0] ? px_buffer_502_r : _GEN_1141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1143 = 10'h1f7 == io_x[9:0] ? px_buffer_503_r : _GEN_1142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1144 = 10'h1f8 == io_x[9:0] ? px_buffer_504_r : _GEN_1143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1145 = 10'h1f9 == io_x[9:0] ? px_buffer_505_r : _GEN_1144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1146 = 10'h1fa == io_x[9:0] ? px_buffer_506_r : _GEN_1145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1147 = 10'h1fb == io_x[9:0] ? px_buffer_507_r : _GEN_1146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1148 = 10'h1fc == io_x[9:0] ? px_buffer_508_r : _GEN_1147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1149 = 10'h1fd == io_x[9:0] ? px_buffer_509_r : _GEN_1148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1150 = 10'h1fe == io_x[9:0] ? px_buffer_510_r : _GEN_1149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1151 = 10'h1ff == io_x[9:0] ? px_buffer_511_r : _GEN_1150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1152 = 10'h200 == io_x[9:0] ? px_buffer_512_r : _GEN_1151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1153 = 10'h201 == io_x[9:0] ? px_buffer_513_r : _GEN_1152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1154 = 10'h202 == io_x[9:0] ? px_buffer_514_r : _GEN_1153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1155 = 10'h203 == io_x[9:0] ? px_buffer_515_r : _GEN_1154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1156 = 10'h204 == io_x[9:0] ? px_buffer_516_r : _GEN_1155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1157 = 10'h205 == io_x[9:0] ? px_buffer_517_r : _GEN_1156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1158 = 10'h206 == io_x[9:0] ? px_buffer_518_r : _GEN_1157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1159 = 10'h207 == io_x[9:0] ? px_buffer_519_r : _GEN_1158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1160 = 10'h208 == io_x[9:0] ? px_buffer_520_r : _GEN_1159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1161 = 10'h209 == io_x[9:0] ? px_buffer_521_r : _GEN_1160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1162 = 10'h20a == io_x[9:0] ? px_buffer_522_r : _GEN_1161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1163 = 10'h20b == io_x[9:0] ? px_buffer_523_r : _GEN_1162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1164 = 10'h20c == io_x[9:0] ? px_buffer_524_r : _GEN_1163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1165 = 10'h20d == io_x[9:0] ? px_buffer_525_r : _GEN_1164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1166 = 10'h20e == io_x[9:0] ? px_buffer_526_r : _GEN_1165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1167 = 10'h20f == io_x[9:0] ? px_buffer_527_r : _GEN_1166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1168 = 10'h210 == io_x[9:0] ? px_buffer_528_r : _GEN_1167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1169 = 10'h211 == io_x[9:0] ? px_buffer_529_r : _GEN_1168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1170 = 10'h212 == io_x[9:0] ? px_buffer_530_r : _GEN_1169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1171 = 10'h213 == io_x[9:0] ? px_buffer_531_r : _GEN_1170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1172 = 10'h214 == io_x[9:0] ? px_buffer_532_r : _GEN_1171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1173 = 10'h215 == io_x[9:0] ? px_buffer_533_r : _GEN_1172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1174 = 10'h216 == io_x[9:0] ? px_buffer_534_r : _GEN_1173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1175 = 10'h217 == io_x[9:0] ? px_buffer_535_r : _GEN_1174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1176 = 10'h218 == io_x[9:0] ? px_buffer_536_r : _GEN_1175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1177 = 10'h219 == io_x[9:0] ? px_buffer_537_r : _GEN_1176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1178 = 10'h21a == io_x[9:0] ? px_buffer_538_r : _GEN_1177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1179 = 10'h21b == io_x[9:0] ? px_buffer_539_r : _GEN_1178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1180 = 10'h21c == io_x[9:0] ? px_buffer_540_r : _GEN_1179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1181 = 10'h21d == io_x[9:0] ? px_buffer_541_r : _GEN_1180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1182 = 10'h21e == io_x[9:0] ? px_buffer_542_r : _GEN_1181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1183 = 10'h21f == io_x[9:0] ? px_buffer_543_r : _GEN_1182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1184 = 10'h220 == io_x[9:0] ? px_buffer_544_r : _GEN_1183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1185 = 10'h221 == io_x[9:0] ? px_buffer_545_r : _GEN_1184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1186 = 10'h222 == io_x[9:0] ? px_buffer_546_r : _GEN_1185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1187 = 10'h223 == io_x[9:0] ? px_buffer_547_r : _GEN_1186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1188 = 10'h224 == io_x[9:0] ? px_buffer_548_r : _GEN_1187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1189 = 10'h225 == io_x[9:0] ? px_buffer_549_r : _GEN_1188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1190 = 10'h226 == io_x[9:0] ? px_buffer_550_r : _GEN_1189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1191 = 10'h227 == io_x[9:0] ? px_buffer_551_r : _GEN_1190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1192 = 10'h228 == io_x[9:0] ? px_buffer_552_r : _GEN_1191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1193 = 10'h229 == io_x[9:0] ? px_buffer_553_r : _GEN_1192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1194 = 10'h22a == io_x[9:0] ? px_buffer_554_r : _GEN_1193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1195 = 10'h22b == io_x[9:0] ? px_buffer_555_r : _GEN_1194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1196 = 10'h22c == io_x[9:0] ? px_buffer_556_r : _GEN_1195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1197 = 10'h22d == io_x[9:0] ? px_buffer_557_r : _GEN_1196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1198 = 10'h22e == io_x[9:0] ? px_buffer_558_r : _GEN_1197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1199 = 10'h22f == io_x[9:0] ? px_buffer_559_r : _GEN_1198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1200 = 10'h230 == io_x[9:0] ? px_buffer_560_r : _GEN_1199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1201 = 10'h231 == io_x[9:0] ? px_buffer_561_r : _GEN_1200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1202 = 10'h232 == io_x[9:0] ? px_buffer_562_r : _GEN_1201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1203 = 10'h233 == io_x[9:0] ? px_buffer_563_r : _GEN_1202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1204 = 10'h234 == io_x[9:0] ? px_buffer_564_r : _GEN_1203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1205 = 10'h235 == io_x[9:0] ? px_buffer_565_r : _GEN_1204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1206 = 10'h236 == io_x[9:0] ? px_buffer_566_r : _GEN_1205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1207 = 10'h237 == io_x[9:0] ? px_buffer_567_r : _GEN_1206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1208 = 10'h238 == io_x[9:0] ? px_buffer_568_r : _GEN_1207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1209 = 10'h239 == io_x[9:0] ? px_buffer_569_r : _GEN_1208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1210 = 10'h23a == io_x[9:0] ? px_buffer_570_r : _GEN_1209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1211 = 10'h23b == io_x[9:0] ? px_buffer_571_r : _GEN_1210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1212 = 10'h23c == io_x[9:0] ? px_buffer_572_r : _GEN_1211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1213 = 10'h23d == io_x[9:0] ? px_buffer_573_r : _GEN_1212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1214 = 10'h23e == io_x[9:0] ? px_buffer_574_r : _GEN_1213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1215 = 10'h23f == io_x[9:0] ? px_buffer_575_r : _GEN_1214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1216 = 10'h240 == io_x[9:0] ? px_buffer_576_r : _GEN_1215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1217 = 10'h241 == io_x[9:0] ? px_buffer_577_r : _GEN_1216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1218 = 10'h242 == io_x[9:0] ? px_buffer_578_r : _GEN_1217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1219 = 10'h243 == io_x[9:0] ? px_buffer_579_r : _GEN_1218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1220 = 10'h244 == io_x[9:0] ? px_buffer_580_r : _GEN_1219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1221 = 10'h245 == io_x[9:0] ? px_buffer_581_r : _GEN_1220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1222 = 10'h246 == io_x[9:0] ? px_buffer_582_r : _GEN_1221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1223 = 10'h247 == io_x[9:0] ? px_buffer_583_r : _GEN_1222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1224 = 10'h248 == io_x[9:0] ? px_buffer_584_r : _GEN_1223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1225 = 10'h249 == io_x[9:0] ? px_buffer_585_r : _GEN_1224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1226 = 10'h24a == io_x[9:0] ? px_buffer_586_r : _GEN_1225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1227 = 10'h24b == io_x[9:0] ? px_buffer_587_r : _GEN_1226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1228 = 10'h24c == io_x[9:0] ? px_buffer_588_r : _GEN_1227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1229 = 10'h24d == io_x[9:0] ? px_buffer_589_r : _GEN_1228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1230 = 10'h24e == io_x[9:0] ? px_buffer_590_r : _GEN_1229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1231 = 10'h24f == io_x[9:0] ? px_buffer_591_r : _GEN_1230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1232 = 10'h250 == io_x[9:0] ? px_buffer_592_r : _GEN_1231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1233 = 10'h251 == io_x[9:0] ? px_buffer_593_r : _GEN_1232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1234 = 10'h252 == io_x[9:0] ? px_buffer_594_r : _GEN_1233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1235 = 10'h253 == io_x[9:0] ? px_buffer_595_r : _GEN_1234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1236 = 10'h254 == io_x[9:0] ? px_buffer_596_r : _GEN_1235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1237 = 10'h255 == io_x[9:0] ? px_buffer_597_r : _GEN_1236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1238 = 10'h256 == io_x[9:0] ? px_buffer_598_r : _GEN_1237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1239 = 10'h257 == io_x[9:0] ? px_buffer_599_r : _GEN_1238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1240 = 10'h258 == io_x[9:0] ? px_buffer_600_r : _GEN_1239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1241 = 10'h259 == io_x[9:0] ? px_buffer_601_r : _GEN_1240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1242 = 10'h25a == io_x[9:0] ? px_buffer_602_r : _GEN_1241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1243 = 10'h25b == io_x[9:0] ? px_buffer_603_r : _GEN_1242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1244 = 10'h25c == io_x[9:0] ? px_buffer_604_r : _GEN_1243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1245 = 10'h25d == io_x[9:0] ? px_buffer_605_r : _GEN_1244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1246 = 10'h25e == io_x[9:0] ? px_buffer_606_r : _GEN_1245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1247 = 10'h25f == io_x[9:0] ? px_buffer_607_r : _GEN_1246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1248 = 10'h260 == io_x[9:0] ? px_buffer_608_r : _GEN_1247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1249 = 10'h261 == io_x[9:0] ? px_buffer_609_r : _GEN_1248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1250 = 10'h262 == io_x[9:0] ? px_buffer_610_r : _GEN_1249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1251 = 10'h263 == io_x[9:0] ? px_buffer_611_r : _GEN_1250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1252 = 10'h264 == io_x[9:0] ? px_buffer_612_r : _GEN_1251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1253 = 10'h265 == io_x[9:0] ? px_buffer_613_r : _GEN_1252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1254 = 10'h266 == io_x[9:0] ? px_buffer_614_r : _GEN_1253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1255 = 10'h267 == io_x[9:0] ? px_buffer_615_r : _GEN_1254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1256 = 10'h268 == io_x[9:0] ? px_buffer_616_r : _GEN_1255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1257 = 10'h269 == io_x[9:0] ? px_buffer_617_r : _GEN_1256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1258 = 10'h26a == io_x[9:0] ? px_buffer_618_r : _GEN_1257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1259 = 10'h26b == io_x[9:0] ? px_buffer_619_r : _GEN_1258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1260 = 10'h26c == io_x[9:0] ? px_buffer_620_r : _GEN_1259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1261 = 10'h26d == io_x[9:0] ? px_buffer_621_r : _GEN_1260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1262 = 10'h26e == io_x[9:0] ? px_buffer_622_r : _GEN_1261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1263 = 10'h26f == io_x[9:0] ? px_buffer_623_r : _GEN_1262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1264 = 10'h270 == io_x[9:0] ? px_buffer_624_r : _GEN_1263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1265 = 10'h271 == io_x[9:0] ? px_buffer_625_r : _GEN_1264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1266 = 10'h272 == io_x[9:0] ? px_buffer_626_r : _GEN_1265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1267 = 10'h273 == io_x[9:0] ? px_buffer_627_r : _GEN_1266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1268 = 10'h274 == io_x[9:0] ? px_buffer_628_r : _GEN_1267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1269 = 10'h275 == io_x[9:0] ? px_buffer_629_r : _GEN_1268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1270 = 10'h276 == io_x[9:0] ? px_buffer_630_r : _GEN_1269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1271 = 10'h277 == io_x[9:0] ? px_buffer_631_r : _GEN_1270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1272 = 10'h278 == io_x[9:0] ? px_buffer_632_r : _GEN_1271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1273 = 10'h279 == io_x[9:0] ? px_buffer_633_r : _GEN_1272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1274 = 10'h27a == io_x[9:0] ? px_buffer_634_r : _GEN_1273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1275 = 10'h27b == io_x[9:0] ? px_buffer_635_r : _GEN_1274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1276 = 10'h27c == io_x[9:0] ? px_buffer_636_r : _GEN_1275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1277 = 10'h27d == io_x[9:0] ? px_buffer_637_r : _GEN_1276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1278 = 10'h27e == io_x[9:0] ? px_buffer_638_r : _GEN_1277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1279 = 10'h27f == io_x[9:0] ? px_buffer_639_r : _GEN_1278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _T_65 = {1'h0,_GEN_1279}; // @[EdgeDetect.scala 55:47]
  wire [8:0] _T_67 = {1'h0,last_px_r}; // @[EdgeDetect.scala 55:79]
  wire [8:0] _T_70 = $signed(_T_65) - $signed(_T_67); // @[EdgeDetect.scala 55:54]
  wire [7:0] _GEN_1281 = 10'h1 == _T_54[9:0] ? px_buffer_1_g : px_buffer_0_g; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1282 = 10'h2 == _T_54[9:0] ? px_buffer_2_g : _GEN_1281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1283 = 10'h3 == _T_54[9:0] ? px_buffer_3_g : _GEN_1282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1284 = 10'h4 == _T_54[9:0] ? px_buffer_4_g : _GEN_1283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1285 = 10'h5 == _T_54[9:0] ? px_buffer_5_g : _GEN_1284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1286 = 10'h6 == _T_54[9:0] ? px_buffer_6_g : _GEN_1285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1287 = 10'h7 == _T_54[9:0] ? px_buffer_7_g : _GEN_1286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1288 = 10'h8 == _T_54[9:0] ? px_buffer_8_g : _GEN_1287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1289 = 10'h9 == _T_54[9:0] ? px_buffer_9_g : _GEN_1288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1290 = 10'ha == _T_54[9:0] ? px_buffer_10_g : _GEN_1289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1291 = 10'hb == _T_54[9:0] ? px_buffer_11_g : _GEN_1290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1292 = 10'hc == _T_54[9:0] ? px_buffer_12_g : _GEN_1291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1293 = 10'hd == _T_54[9:0] ? px_buffer_13_g : _GEN_1292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1294 = 10'he == _T_54[9:0] ? px_buffer_14_g : _GEN_1293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1295 = 10'hf == _T_54[9:0] ? px_buffer_15_g : _GEN_1294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1296 = 10'h10 == _T_54[9:0] ? px_buffer_16_g : _GEN_1295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1297 = 10'h11 == _T_54[9:0] ? px_buffer_17_g : _GEN_1296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1298 = 10'h12 == _T_54[9:0] ? px_buffer_18_g : _GEN_1297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1299 = 10'h13 == _T_54[9:0] ? px_buffer_19_g : _GEN_1298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1300 = 10'h14 == _T_54[9:0] ? px_buffer_20_g : _GEN_1299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1301 = 10'h15 == _T_54[9:0] ? px_buffer_21_g : _GEN_1300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1302 = 10'h16 == _T_54[9:0] ? px_buffer_22_g : _GEN_1301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1303 = 10'h17 == _T_54[9:0] ? px_buffer_23_g : _GEN_1302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1304 = 10'h18 == _T_54[9:0] ? px_buffer_24_g : _GEN_1303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1305 = 10'h19 == _T_54[9:0] ? px_buffer_25_g : _GEN_1304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1306 = 10'h1a == _T_54[9:0] ? px_buffer_26_g : _GEN_1305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1307 = 10'h1b == _T_54[9:0] ? px_buffer_27_g : _GEN_1306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1308 = 10'h1c == _T_54[9:0] ? px_buffer_28_g : _GEN_1307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1309 = 10'h1d == _T_54[9:0] ? px_buffer_29_g : _GEN_1308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1310 = 10'h1e == _T_54[9:0] ? px_buffer_30_g : _GEN_1309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1311 = 10'h1f == _T_54[9:0] ? px_buffer_31_g : _GEN_1310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1312 = 10'h20 == _T_54[9:0] ? px_buffer_32_g : _GEN_1311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1313 = 10'h21 == _T_54[9:0] ? px_buffer_33_g : _GEN_1312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1314 = 10'h22 == _T_54[9:0] ? px_buffer_34_g : _GEN_1313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1315 = 10'h23 == _T_54[9:0] ? px_buffer_35_g : _GEN_1314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1316 = 10'h24 == _T_54[9:0] ? px_buffer_36_g : _GEN_1315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1317 = 10'h25 == _T_54[9:0] ? px_buffer_37_g : _GEN_1316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1318 = 10'h26 == _T_54[9:0] ? px_buffer_38_g : _GEN_1317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1319 = 10'h27 == _T_54[9:0] ? px_buffer_39_g : _GEN_1318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1320 = 10'h28 == _T_54[9:0] ? px_buffer_40_g : _GEN_1319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1321 = 10'h29 == _T_54[9:0] ? px_buffer_41_g : _GEN_1320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1322 = 10'h2a == _T_54[9:0] ? px_buffer_42_g : _GEN_1321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1323 = 10'h2b == _T_54[9:0] ? px_buffer_43_g : _GEN_1322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1324 = 10'h2c == _T_54[9:0] ? px_buffer_44_g : _GEN_1323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1325 = 10'h2d == _T_54[9:0] ? px_buffer_45_g : _GEN_1324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1326 = 10'h2e == _T_54[9:0] ? px_buffer_46_g : _GEN_1325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1327 = 10'h2f == _T_54[9:0] ? px_buffer_47_g : _GEN_1326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1328 = 10'h30 == _T_54[9:0] ? px_buffer_48_g : _GEN_1327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1329 = 10'h31 == _T_54[9:0] ? px_buffer_49_g : _GEN_1328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1330 = 10'h32 == _T_54[9:0] ? px_buffer_50_g : _GEN_1329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1331 = 10'h33 == _T_54[9:0] ? px_buffer_51_g : _GEN_1330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1332 = 10'h34 == _T_54[9:0] ? px_buffer_52_g : _GEN_1331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1333 = 10'h35 == _T_54[9:0] ? px_buffer_53_g : _GEN_1332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1334 = 10'h36 == _T_54[9:0] ? px_buffer_54_g : _GEN_1333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1335 = 10'h37 == _T_54[9:0] ? px_buffer_55_g : _GEN_1334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1336 = 10'h38 == _T_54[9:0] ? px_buffer_56_g : _GEN_1335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1337 = 10'h39 == _T_54[9:0] ? px_buffer_57_g : _GEN_1336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1338 = 10'h3a == _T_54[9:0] ? px_buffer_58_g : _GEN_1337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1339 = 10'h3b == _T_54[9:0] ? px_buffer_59_g : _GEN_1338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1340 = 10'h3c == _T_54[9:0] ? px_buffer_60_g : _GEN_1339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1341 = 10'h3d == _T_54[9:0] ? px_buffer_61_g : _GEN_1340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1342 = 10'h3e == _T_54[9:0] ? px_buffer_62_g : _GEN_1341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1343 = 10'h3f == _T_54[9:0] ? px_buffer_63_g : _GEN_1342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1344 = 10'h40 == _T_54[9:0] ? px_buffer_64_g : _GEN_1343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1345 = 10'h41 == _T_54[9:0] ? px_buffer_65_g : _GEN_1344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1346 = 10'h42 == _T_54[9:0] ? px_buffer_66_g : _GEN_1345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1347 = 10'h43 == _T_54[9:0] ? px_buffer_67_g : _GEN_1346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1348 = 10'h44 == _T_54[9:0] ? px_buffer_68_g : _GEN_1347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1349 = 10'h45 == _T_54[9:0] ? px_buffer_69_g : _GEN_1348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1350 = 10'h46 == _T_54[9:0] ? px_buffer_70_g : _GEN_1349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1351 = 10'h47 == _T_54[9:0] ? px_buffer_71_g : _GEN_1350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1352 = 10'h48 == _T_54[9:0] ? px_buffer_72_g : _GEN_1351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1353 = 10'h49 == _T_54[9:0] ? px_buffer_73_g : _GEN_1352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1354 = 10'h4a == _T_54[9:0] ? px_buffer_74_g : _GEN_1353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1355 = 10'h4b == _T_54[9:0] ? px_buffer_75_g : _GEN_1354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1356 = 10'h4c == _T_54[9:0] ? px_buffer_76_g : _GEN_1355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1357 = 10'h4d == _T_54[9:0] ? px_buffer_77_g : _GEN_1356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1358 = 10'h4e == _T_54[9:0] ? px_buffer_78_g : _GEN_1357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1359 = 10'h4f == _T_54[9:0] ? px_buffer_79_g : _GEN_1358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1360 = 10'h50 == _T_54[9:0] ? px_buffer_80_g : _GEN_1359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1361 = 10'h51 == _T_54[9:0] ? px_buffer_81_g : _GEN_1360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1362 = 10'h52 == _T_54[9:0] ? px_buffer_82_g : _GEN_1361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1363 = 10'h53 == _T_54[9:0] ? px_buffer_83_g : _GEN_1362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1364 = 10'h54 == _T_54[9:0] ? px_buffer_84_g : _GEN_1363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1365 = 10'h55 == _T_54[9:0] ? px_buffer_85_g : _GEN_1364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1366 = 10'h56 == _T_54[9:0] ? px_buffer_86_g : _GEN_1365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1367 = 10'h57 == _T_54[9:0] ? px_buffer_87_g : _GEN_1366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1368 = 10'h58 == _T_54[9:0] ? px_buffer_88_g : _GEN_1367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1369 = 10'h59 == _T_54[9:0] ? px_buffer_89_g : _GEN_1368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1370 = 10'h5a == _T_54[9:0] ? px_buffer_90_g : _GEN_1369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1371 = 10'h5b == _T_54[9:0] ? px_buffer_91_g : _GEN_1370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1372 = 10'h5c == _T_54[9:0] ? px_buffer_92_g : _GEN_1371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1373 = 10'h5d == _T_54[9:0] ? px_buffer_93_g : _GEN_1372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1374 = 10'h5e == _T_54[9:0] ? px_buffer_94_g : _GEN_1373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1375 = 10'h5f == _T_54[9:0] ? px_buffer_95_g : _GEN_1374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1376 = 10'h60 == _T_54[9:0] ? px_buffer_96_g : _GEN_1375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1377 = 10'h61 == _T_54[9:0] ? px_buffer_97_g : _GEN_1376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1378 = 10'h62 == _T_54[9:0] ? px_buffer_98_g : _GEN_1377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1379 = 10'h63 == _T_54[9:0] ? px_buffer_99_g : _GEN_1378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1380 = 10'h64 == _T_54[9:0] ? px_buffer_100_g : _GEN_1379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1381 = 10'h65 == _T_54[9:0] ? px_buffer_101_g : _GEN_1380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1382 = 10'h66 == _T_54[9:0] ? px_buffer_102_g : _GEN_1381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1383 = 10'h67 == _T_54[9:0] ? px_buffer_103_g : _GEN_1382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1384 = 10'h68 == _T_54[9:0] ? px_buffer_104_g : _GEN_1383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1385 = 10'h69 == _T_54[9:0] ? px_buffer_105_g : _GEN_1384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1386 = 10'h6a == _T_54[9:0] ? px_buffer_106_g : _GEN_1385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1387 = 10'h6b == _T_54[9:0] ? px_buffer_107_g : _GEN_1386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1388 = 10'h6c == _T_54[9:0] ? px_buffer_108_g : _GEN_1387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1389 = 10'h6d == _T_54[9:0] ? px_buffer_109_g : _GEN_1388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1390 = 10'h6e == _T_54[9:0] ? px_buffer_110_g : _GEN_1389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1391 = 10'h6f == _T_54[9:0] ? px_buffer_111_g : _GEN_1390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1392 = 10'h70 == _T_54[9:0] ? px_buffer_112_g : _GEN_1391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1393 = 10'h71 == _T_54[9:0] ? px_buffer_113_g : _GEN_1392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1394 = 10'h72 == _T_54[9:0] ? px_buffer_114_g : _GEN_1393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1395 = 10'h73 == _T_54[9:0] ? px_buffer_115_g : _GEN_1394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1396 = 10'h74 == _T_54[9:0] ? px_buffer_116_g : _GEN_1395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1397 = 10'h75 == _T_54[9:0] ? px_buffer_117_g : _GEN_1396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1398 = 10'h76 == _T_54[9:0] ? px_buffer_118_g : _GEN_1397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1399 = 10'h77 == _T_54[9:0] ? px_buffer_119_g : _GEN_1398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1400 = 10'h78 == _T_54[9:0] ? px_buffer_120_g : _GEN_1399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1401 = 10'h79 == _T_54[9:0] ? px_buffer_121_g : _GEN_1400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1402 = 10'h7a == _T_54[9:0] ? px_buffer_122_g : _GEN_1401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1403 = 10'h7b == _T_54[9:0] ? px_buffer_123_g : _GEN_1402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1404 = 10'h7c == _T_54[9:0] ? px_buffer_124_g : _GEN_1403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1405 = 10'h7d == _T_54[9:0] ? px_buffer_125_g : _GEN_1404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1406 = 10'h7e == _T_54[9:0] ? px_buffer_126_g : _GEN_1405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1407 = 10'h7f == _T_54[9:0] ? px_buffer_127_g : _GEN_1406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1408 = 10'h80 == _T_54[9:0] ? px_buffer_128_g : _GEN_1407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1409 = 10'h81 == _T_54[9:0] ? px_buffer_129_g : _GEN_1408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1410 = 10'h82 == _T_54[9:0] ? px_buffer_130_g : _GEN_1409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1411 = 10'h83 == _T_54[9:0] ? px_buffer_131_g : _GEN_1410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1412 = 10'h84 == _T_54[9:0] ? px_buffer_132_g : _GEN_1411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1413 = 10'h85 == _T_54[9:0] ? px_buffer_133_g : _GEN_1412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1414 = 10'h86 == _T_54[9:0] ? px_buffer_134_g : _GEN_1413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1415 = 10'h87 == _T_54[9:0] ? px_buffer_135_g : _GEN_1414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1416 = 10'h88 == _T_54[9:0] ? px_buffer_136_g : _GEN_1415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1417 = 10'h89 == _T_54[9:0] ? px_buffer_137_g : _GEN_1416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1418 = 10'h8a == _T_54[9:0] ? px_buffer_138_g : _GEN_1417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1419 = 10'h8b == _T_54[9:0] ? px_buffer_139_g : _GEN_1418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1420 = 10'h8c == _T_54[9:0] ? px_buffer_140_g : _GEN_1419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1421 = 10'h8d == _T_54[9:0] ? px_buffer_141_g : _GEN_1420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1422 = 10'h8e == _T_54[9:0] ? px_buffer_142_g : _GEN_1421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1423 = 10'h8f == _T_54[9:0] ? px_buffer_143_g : _GEN_1422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1424 = 10'h90 == _T_54[9:0] ? px_buffer_144_g : _GEN_1423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1425 = 10'h91 == _T_54[9:0] ? px_buffer_145_g : _GEN_1424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1426 = 10'h92 == _T_54[9:0] ? px_buffer_146_g : _GEN_1425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1427 = 10'h93 == _T_54[9:0] ? px_buffer_147_g : _GEN_1426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1428 = 10'h94 == _T_54[9:0] ? px_buffer_148_g : _GEN_1427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1429 = 10'h95 == _T_54[9:0] ? px_buffer_149_g : _GEN_1428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1430 = 10'h96 == _T_54[9:0] ? px_buffer_150_g : _GEN_1429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1431 = 10'h97 == _T_54[9:0] ? px_buffer_151_g : _GEN_1430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1432 = 10'h98 == _T_54[9:0] ? px_buffer_152_g : _GEN_1431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1433 = 10'h99 == _T_54[9:0] ? px_buffer_153_g : _GEN_1432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1434 = 10'h9a == _T_54[9:0] ? px_buffer_154_g : _GEN_1433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1435 = 10'h9b == _T_54[9:0] ? px_buffer_155_g : _GEN_1434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1436 = 10'h9c == _T_54[9:0] ? px_buffer_156_g : _GEN_1435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1437 = 10'h9d == _T_54[9:0] ? px_buffer_157_g : _GEN_1436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1438 = 10'h9e == _T_54[9:0] ? px_buffer_158_g : _GEN_1437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1439 = 10'h9f == _T_54[9:0] ? px_buffer_159_g : _GEN_1438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1440 = 10'ha0 == _T_54[9:0] ? px_buffer_160_g : _GEN_1439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1441 = 10'ha1 == _T_54[9:0] ? px_buffer_161_g : _GEN_1440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1442 = 10'ha2 == _T_54[9:0] ? px_buffer_162_g : _GEN_1441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1443 = 10'ha3 == _T_54[9:0] ? px_buffer_163_g : _GEN_1442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1444 = 10'ha4 == _T_54[9:0] ? px_buffer_164_g : _GEN_1443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1445 = 10'ha5 == _T_54[9:0] ? px_buffer_165_g : _GEN_1444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1446 = 10'ha6 == _T_54[9:0] ? px_buffer_166_g : _GEN_1445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1447 = 10'ha7 == _T_54[9:0] ? px_buffer_167_g : _GEN_1446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1448 = 10'ha8 == _T_54[9:0] ? px_buffer_168_g : _GEN_1447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1449 = 10'ha9 == _T_54[9:0] ? px_buffer_169_g : _GEN_1448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1450 = 10'haa == _T_54[9:0] ? px_buffer_170_g : _GEN_1449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1451 = 10'hab == _T_54[9:0] ? px_buffer_171_g : _GEN_1450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1452 = 10'hac == _T_54[9:0] ? px_buffer_172_g : _GEN_1451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1453 = 10'had == _T_54[9:0] ? px_buffer_173_g : _GEN_1452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1454 = 10'hae == _T_54[9:0] ? px_buffer_174_g : _GEN_1453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1455 = 10'haf == _T_54[9:0] ? px_buffer_175_g : _GEN_1454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1456 = 10'hb0 == _T_54[9:0] ? px_buffer_176_g : _GEN_1455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1457 = 10'hb1 == _T_54[9:0] ? px_buffer_177_g : _GEN_1456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1458 = 10'hb2 == _T_54[9:0] ? px_buffer_178_g : _GEN_1457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1459 = 10'hb3 == _T_54[9:0] ? px_buffer_179_g : _GEN_1458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1460 = 10'hb4 == _T_54[9:0] ? px_buffer_180_g : _GEN_1459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1461 = 10'hb5 == _T_54[9:0] ? px_buffer_181_g : _GEN_1460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1462 = 10'hb6 == _T_54[9:0] ? px_buffer_182_g : _GEN_1461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1463 = 10'hb7 == _T_54[9:0] ? px_buffer_183_g : _GEN_1462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1464 = 10'hb8 == _T_54[9:0] ? px_buffer_184_g : _GEN_1463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1465 = 10'hb9 == _T_54[9:0] ? px_buffer_185_g : _GEN_1464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1466 = 10'hba == _T_54[9:0] ? px_buffer_186_g : _GEN_1465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1467 = 10'hbb == _T_54[9:0] ? px_buffer_187_g : _GEN_1466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1468 = 10'hbc == _T_54[9:0] ? px_buffer_188_g : _GEN_1467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1469 = 10'hbd == _T_54[9:0] ? px_buffer_189_g : _GEN_1468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1470 = 10'hbe == _T_54[9:0] ? px_buffer_190_g : _GEN_1469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1471 = 10'hbf == _T_54[9:0] ? px_buffer_191_g : _GEN_1470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1472 = 10'hc0 == _T_54[9:0] ? px_buffer_192_g : _GEN_1471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1473 = 10'hc1 == _T_54[9:0] ? px_buffer_193_g : _GEN_1472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1474 = 10'hc2 == _T_54[9:0] ? px_buffer_194_g : _GEN_1473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1475 = 10'hc3 == _T_54[9:0] ? px_buffer_195_g : _GEN_1474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1476 = 10'hc4 == _T_54[9:0] ? px_buffer_196_g : _GEN_1475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1477 = 10'hc5 == _T_54[9:0] ? px_buffer_197_g : _GEN_1476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1478 = 10'hc6 == _T_54[9:0] ? px_buffer_198_g : _GEN_1477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1479 = 10'hc7 == _T_54[9:0] ? px_buffer_199_g : _GEN_1478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1480 = 10'hc8 == _T_54[9:0] ? px_buffer_200_g : _GEN_1479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1481 = 10'hc9 == _T_54[9:0] ? px_buffer_201_g : _GEN_1480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1482 = 10'hca == _T_54[9:0] ? px_buffer_202_g : _GEN_1481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1483 = 10'hcb == _T_54[9:0] ? px_buffer_203_g : _GEN_1482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1484 = 10'hcc == _T_54[9:0] ? px_buffer_204_g : _GEN_1483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1485 = 10'hcd == _T_54[9:0] ? px_buffer_205_g : _GEN_1484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1486 = 10'hce == _T_54[9:0] ? px_buffer_206_g : _GEN_1485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1487 = 10'hcf == _T_54[9:0] ? px_buffer_207_g : _GEN_1486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1488 = 10'hd0 == _T_54[9:0] ? px_buffer_208_g : _GEN_1487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1489 = 10'hd1 == _T_54[9:0] ? px_buffer_209_g : _GEN_1488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1490 = 10'hd2 == _T_54[9:0] ? px_buffer_210_g : _GEN_1489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1491 = 10'hd3 == _T_54[9:0] ? px_buffer_211_g : _GEN_1490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1492 = 10'hd4 == _T_54[9:0] ? px_buffer_212_g : _GEN_1491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1493 = 10'hd5 == _T_54[9:0] ? px_buffer_213_g : _GEN_1492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1494 = 10'hd6 == _T_54[9:0] ? px_buffer_214_g : _GEN_1493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1495 = 10'hd7 == _T_54[9:0] ? px_buffer_215_g : _GEN_1494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1496 = 10'hd8 == _T_54[9:0] ? px_buffer_216_g : _GEN_1495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1497 = 10'hd9 == _T_54[9:0] ? px_buffer_217_g : _GEN_1496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1498 = 10'hda == _T_54[9:0] ? px_buffer_218_g : _GEN_1497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1499 = 10'hdb == _T_54[9:0] ? px_buffer_219_g : _GEN_1498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1500 = 10'hdc == _T_54[9:0] ? px_buffer_220_g : _GEN_1499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1501 = 10'hdd == _T_54[9:0] ? px_buffer_221_g : _GEN_1500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1502 = 10'hde == _T_54[9:0] ? px_buffer_222_g : _GEN_1501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1503 = 10'hdf == _T_54[9:0] ? px_buffer_223_g : _GEN_1502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1504 = 10'he0 == _T_54[9:0] ? px_buffer_224_g : _GEN_1503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1505 = 10'he1 == _T_54[9:0] ? px_buffer_225_g : _GEN_1504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1506 = 10'he2 == _T_54[9:0] ? px_buffer_226_g : _GEN_1505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1507 = 10'he3 == _T_54[9:0] ? px_buffer_227_g : _GEN_1506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1508 = 10'he4 == _T_54[9:0] ? px_buffer_228_g : _GEN_1507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1509 = 10'he5 == _T_54[9:0] ? px_buffer_229_g : _GEN_1508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1510 = 10'he6 == _T_54[9:0] ? px_buffer_230_g : _GEN_1509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1511 = 10'he7 == _T_54[9:0] ? px_buffer_231_g : _GEN_1510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1512 = 10'he8 == _T_54[9:0] ? px_buffer_232_g : _GEN_1511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1513 = 10'he9 == _T_54[9:0] ? px_buffer_233_g : _GEN_1512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1514 = 10'hea == _T_54[9:0] ? px_buffer_234_g : _GEN_1513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1515 = 10'heb == _T_54[9:0] ? px_buffer_235_g : _GEN_1514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1516 = 10'hec == _T_54[9:0] ? px_buffer_236_g : _GEN_1515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1517 = 10'hed == _T_54[9:0] ? px_buffer_237_g : _GEN_1516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1518 = 10'hee == _T_54[9:0] ? px_buffer_238_g : _GEN_1517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1519 = 10'hef == _T_54[9:0] ? px_buffer_239_g : _GEN_1518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1520 = 10'hf0 == _T_54[9:0] ? px_buffer_240_g : _GEN_1519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1521 = 10'hf1 == _T_54[9:0] ? px_buffer_241_g : _GEN_1520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1522 = 10'hf2 == _T_54[9:0] ? px_buffer_242_g : _GEN_1521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1523 = 10'hf3 == _T_54[9:0] ? px_buffer_243_g : _GEN_1522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1524 = 10'hf4 == _T_54[9:0] ? px_buffer_244_g : _GEN_1523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1525 = 10'hf5 == _T_54[9:0] ? px_buffer_245_g : _GEN_1524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1526 = 10'hf6 == _T_54[9:0] ? px_buffer_246_g : _GEN_1525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1527 = 10'hf7 == _T_54[9:0] ? px_buffer_247_g : _GEN_1526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1528 = 10'hf8 == _T_54[9:0] ? px_buffer_248_g : _GEN_1527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1529 = 10'hf9 == _T_54[9:0] ? px_buffer_249_g : _GEN_1528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1530 = 10'hfa == _T_54[9:0] ? px_buffer_250_g : _GEN_1529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1531 = 10'hfb == _T_54[9:0] ? px_buffer_251_g : _GEN_1530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1532 = 10'hfc == _T_54[9:0] ? px_buffer_252_g : _GEN_1531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1533 = 10'hfd == _T_54[9:0] ? px_buffer_253_g : _GEN_1532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1534 = 10'hfe == _T_54[9:0] ? px_buffer_254_g : _GEN_1533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1535 = 10'hff == _T_54[9:0] ? px_buffer_255_g : _GEN_1534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1536 = 10'h100 == _T_54[9:0] ? px_buffer_256_g : _GEN_1535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1537 = 10'h101 == _T_54[9:0] ? px_buffer_257_g : _GEN_1536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1538 = 10'h102 == _T_54[9:0] ? px_buffer_258_g : _GEN_1537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1539 = 10'h103 == _T_54[9:0] ? px_buffer_259_g : _GEN_1538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1540 = 10'h104 == _T_54[9:0] ? px_buffer_260_g : _GEN_1539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1541 = 10'h105 == _T_54[9:0] ? px_buffer_261_g : _GEN_1540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1542 = 10'h106 == _T_54[9:0] ? px_buffer_262_g : _GEN_1541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1543 = 10'h107 == _T_54[9:0] ? px_buffer_263_g : _GEN_1542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1544 = 10'h108 == _T_54[9:0] ? px_buffer_264_g : _GEN_1543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1545 = 10'h109 == _T_54[9:0] ? px_buffer_265_g : _GEN_1544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1546 = 10'h10a == _T_54[9:0] ? px_buffer_266_g : _GEN_1545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1547 = 10'h10b == _T_54[9:0] ? px_buffer_267_g : _GEN_1546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1548 = 10'h10c == _T_54[9:0] ? px_buffer_268_g : _GEN_1547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1549 = 10'h10d == _T_54[9:0] ? px_buffer_269_g : _GEN_1548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1550 = 10'h10e == _T_54[9:0] ? px_buffer_270_g : _GEN_1549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1551 = 10'h10f == _T_54[9:0] ? px_buffer_271_g : _GEN_1550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1552 = 10'h110 == _T_54[9:0] ? px_buffer_272_g : _GEN_1551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1553 = 10'h111 == _T_54[9:0] ? px_buffer_273_g : _GEN_1552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1554 = 10'h112 == _T_54[9:0] ? px_buffer_274_g : _GEN_1553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1555 = 10'h113 == _T_54[9:0] ? px_buffer_275_g : _GEN_1554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1556 = 10'h114 == _T_54[9:0] ? px_buffer_276_g : _GEN_1555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1557 = 10'h115 == _T_54[9:0] ? px_buffer_277_g : _GEN_1556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1558 = 10'h116 == _T_54[9:0] ? px_buffer_278_g : _GEN_1557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1559 = 10'h117 == _T_54[9:0] ? px_buffer_279_g : _GEN_1558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1560 = 10'h118 == _T_54[9:0] ? px_buffer_280_g : _GEN_1559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1561 = 10'h119 == _T_54[9:0] ? px_buffer_281_g : _GEN_1560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1562 = 10'h11a == _T_54[9:0] ? px_buffer_282_g : _GEN_1561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1563 = 10'h11b == _T_54[9:0] ? px_buffer_283_g : _GEN_1562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1564 = 10'h11c == _T_54[9:0] ? px_buffer_284_g : _GEN_1563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1565 = 10'h11d == _T_54[9:0] ? px_buffer_285_g : _GEN_1564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1566 = 10'h11e == _T_54[9:0] ? px_buffer_286_g : _GEN_1565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1567 = 10'h11f == _T_54[9:0] ? px_buffer_287_g : _GEN_1566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1568 = 10'h120 == _T_54[9:0] ? px_buffer_288_g : _GEN_1567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1569 = 10'h121 == _T_54[9:0] ? px_buffer_289_g : _GEN_1568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1570 = 10'h122 == _T_54[9:0] ? px_buffer_290_g : _GEN_1569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1571 = 10'h123 == _T_54[9:0] ? px_buffer_291_g : _GEN_1570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1572 = 10'h124 == _T_54[9:0] ? px_buffer_292_g : _GEN_1571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1573 = 10'h125 == _T_54[9:0] ? px_buffer_293_g : _GEN_1572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1574 = 10'h126 == _T_54[9:0] ? px_buffer_294_g : _GEN_1573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1575 = 10'h127 == _T_54[9:0] ? px_buffer_295_g : _GEN_1574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1576 = 10'h128 == _T_54[9:0] ? px_buffer_296_g : _GEN_1575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1577 = 10'h129 == _T_54[9:0] ? px_buffer_297_g : _GEN_1576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1578 = 10'h12a == _T_54[9:0] ? px_buffer_298_g : _GEN_1577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1579 = 10'h12b == _T_54[9:0] ? px_buffer_299_g : _GEN_1578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1580 = 10'h12c == _T_54[9:0] ? px_buffer_300_g : _GEN_1579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1581 = 10'h12d == _T_54[9:0] ? px_buffer_301_g : _GEN_1580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1582 = 10'h12e == _T_54[9:0] ? px_buffer_302_g : _GEN_1581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1583 = 10'h12f == _T_54[9:0] ? px_buffer_303_g : _GEN_1582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1584 = 10'h130 == _T_54[9:0] ? px_buffer_304_g : _GEN_1583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1585 = 10'h131 == _T_54[9:0] ? px_buffer_305_g : _GEN_1584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1586 = 10'h132 == _T_54[9:0] ? px_buffer_306_g : _GEN_1585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1587 = 10'h133 == _T_54[9:0] ? px_buffer_307_g : _GEN_1586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1588 = 10'h134 == _T_54[9:0] ? px_buffer_308_g : _GEN_1587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1589 = 10'h135 == _T_54[9:0] ? px_buffer_309_g : _GEN_1588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1590 = 10'h136 == _T_54[9:0] ? px_buffer_310_g : _GEN_1589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1591 = 10'h137 == _T_54[9:0] ? px_buffer_311_g : _GEN_1590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1592 = 10'h138 == _T_54[9:0] ? px_buffer_312_g : _GEN_1591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1593 = 10'h139 == _T_54[9:0] ? px_buffer_313_g : _GEN_1592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1594 = 10'h13a == _T_54[9:0] ? px_buffer_314_g : _GEN_1593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1595 = 10'h13b == _T_54[9:0] ? px_buffer_315_g : _GEN_1594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1596 = 10'h13c == _T_54[9:0] ? px_buffer_316_g : _GEN_1595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1597 = 10'h13d == _T_54[9:0] ? px_buffer_317_g : _GEN_1596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1598 = 10'h13e == _T_54[9:0] ? px_buffer_318_g : _GEN_1597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1599 = 10'h13f == _T_54[9:0] ? px_buffer_319_g : _GEN_1598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1600 = 10'h140 == _T_54[9:0] ? px_buffer_320_g : _GEN_1599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1601 = 10'h141 == _T_54[9:0] ? px_buffer_321_g : _GEN_1600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1602 = 10'h142 == _T_54[9:0] ? px_buffer_322_g : _GEN_1601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1603 = 10'h143 == _T_54[9:0] ? px_buffer_323_g : _GEN_1602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1604 = 10'h144 == _T_54[9:0] ? px_buffer_324_g : _GEN_1603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1605 = 10'h145 == _T_54[9:0] ? px_buffer_325_g : _GEN_1604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1606 = 10'h146 == _T_54[9:0] ? px_buffer_326_g : _GEN_1605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1607 = 10'h147 == _T_54[9:0] ? px_buffer_327_g : _GEN_1606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1608 = 10'h148 == _T_54[9:0] ? px_buffer_328_g : _GEN_1607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1609 = 10'h149 == _T_54[9:0] ? px_buffer_329_g : _GEN_1608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1610 = 10'h14a == _T_54[9:0] ? px_buffer_330_g : _GEN_1609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1611 = 10'h14b == _T_54[9:0] ? px_buffer_331_g : _GEN_1610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1612 = 10'h14c == _T_54[9:0] ? px_buffer_332_g : _GEN_1611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1613 = 10'h14d == _T_54[9:0] ? px_buffer_333_g : _GEN_1612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1614 = 10'h14e == _T_54[9:0] ? px_buffer_334_g : _GEN_1613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1615 = 10'h14f == _T_54[9:0] ? px_buffer_335_g : _GEN_1614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1616 = 10'h150 == _T_54[9:0] ? px_buffer_336_g : _GEN_1615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1617 = 10'h151 == _T_54[9:0] ? px_buffer_337_g : _GEN_1616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1618 = 10'h152 == _T_54[9:0] ? px_buffer_338_g : _GEN_1617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1619 = 10'h153 == _T_54[9:0] ? px_buffer_339_g : _GEN_1618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1620 = 10'h154 == _T_54[9:0] ? px_buffer_340_g : _GEN_1619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1621 = 10'h155 == _T_54[9:0] ? px_buffer_341_g : _GEN_1620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1622 = 10'h156 == _T_54[9:0] ? px_buffer_342_g : _GEN_1621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1623 = 10'h157 == _T_54[9:0] ? px_buffer_343_g : _GEN_1622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1624 = 10'h158 == _T_54[9:0] ? px_buffer_344_g : _GEN_1623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1625 = 10'h159 == _T_54[9:0] ? px_buffer_345_g : _GEN_1624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1626 = 10'h15a == _T_54[9:0] ? px_buffer_346_g : _GEN_1625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1627 = 10'h15b == _T_54[9:0] ? px_buffer_347_g : _GEN_1626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1628 = 10'h15c == _T_54[9:0] ? px_buffer_348_g : _GEN_1627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1629 = 10'h15d == _T_54[9:0] ? px_buffer_349_g : _GEN_1628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1630 = 10'h15e == _T_54[9:0] ? px_buffer_350_g : _GEN_1629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1631 = 10'h15f == _T_54[9:0] ? px_buffer_351_g : _GEN_1630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1632 = 10'h160 == _T_54[9:0] ? px_buffer_352_g : _GEN_1631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1633 = 10'h161 == _T_54[9:0] ? px_buffer_353_g : _GEN_1632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1634 = 10'h162 == _T_54[9:0] ? px_buffer_354_g : _GEN_1633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1635 = 10'h163 == _T_54[9:0] ? px_buffer_355_g : _GEN_1634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1636 = 10'h164 == _T_54[9:0] ? px_buffer_356_g : _GEN_1635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1637 = 10'h165 == _T_54[9:0] ? px_buffer_357_g : _GEN_1636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1638 = 10'h166 == _T_54[9:0] ? px_buffer_358_g : _GEN_1637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1639 = 10'h167 == _T_54[9:0] ? px_buffer_359_g : _GEN_1638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1640 = 10'h168 == _T_54[9:0] ? px_buffer_360_g : _GEN_1639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1641 = 10'h169 == _T_54[9:0] ? px_buffer_361_g : _GEN_1640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1642 = 10'h16a == _T_54[9:0] ? px_buffer_362_g : _GEN_1641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1643 = 10'h16b == _T_54[9:0] ? px_buffer_363_g : _GEN_1642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1644 = 10'h16c == _T_54[9:0] ? px_buffer_364_g : _GEN_1643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1645 = 10'h16d == _T_54[9:0] ? px_buffer_365_g : _GEN_1644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1646 = 10'h16e == _T_54[9:0] ? px_buffer_366_g : _GEN_1645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1647 = 10'h16f == _T_54[9:0] ? px_buffer_367_g : _GEN_1646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1648 = 10'h170 == _T_54[9:0] ? px_buffer_368_g : _GEN_1647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1649 = 10'h171 == _T_54[9:0] ? px_buffer_369_g : _GEN_1648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1650 = 10'h172 == _T_54[9:0] ? px_buffer_370_g : _GEN_1649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1651 = 10'h173 == _T_54[9:0] ? px_buffer_371_g : _GEN_1650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1652 = 10'h174 == _T_54[9:0] ? px_buffer_372_g : _GEN_1651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1653 = 10'h175 == _T_54[9:0] ? px_buffer_373_g : _GEN_1652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1654 = 10'h176 == _T_54[9:0] ? px_buffer_374_g : _GEN_1653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1655 = 10'h177 == _T_54[9:0] ? px_buffer_375_g : _GEN_1654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1656 = 10'h178 == _T_54[9:0] ? px_buffer_376_g : _GEN_1655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1657 = 10'h179 == _T_54[9:0] ? px_buffer_377_g : _GEN_1656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1658 = 10'h17a == _T_54[9:0] ? px_buffer_378_g : _GEN_1657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1659 = 10'h17b == _T_54[9:0] ? px_buffer_379_g : _GEN_1658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1660 = 10'h17c == _T_54[9:0] ? px_buffer_380_g : _GEN_1659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1661 = 10'h17d == _T_54[9:0] ? px_buffer_381_g : _GEN_1660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1662 = 10'h17e == _T_54[9:0] ? px_buffer_382_g : _GEN_1661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1663 = 10'h17f == _T_54[9:0] ? px_buffer_383_g : _GEN_1662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1664 = 10'h180 == _T_54[9:0] ? px_buffer_384_g : _GEN_1663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1665 = 10'h181 == _T_54[9:0] ? px_buffer_385_g : _GEN_1664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1666 = 10'h182 == _T_54[9:0] ? px_buffer_386_g : _GEN_1665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1667 = 10'h183 == _T_54[9:0] ? px_buffer_387_g : _GEN_1666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1668 = 10'h184 == _T_54[9:0] ? px_buffer_388_g : _GEN_1667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1669 = 10'h185 == _T_54[9:0] ? px_buffer_389_g : _GEN_1668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1670 = 10'h186 == _T_54[9:0] ? px_buffer_390_g : _GEN_1669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1671 = 10'h187 == _T_54[9:0] ? px_buffer_391_g : _GEN_1670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1672 = 10'h188 == _T_54[9:0] ? px_buffer_392_g : _GEN_1671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1673 = 10'h189 == _T_54[9:0] ? px_buffer_393_g : _GEN_1672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1674 = 10'h18a == _T_54[9:0] ? px_buffer_394_g : _GEN_1673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1675 = 10'h18b == _T_54[9:0] ? px_buffer_395_g : _GEN_1674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1676 = 10'h18c == _T_54[9:0] ? px_buffer_396_g : _GEN_1675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1677 = 10'h18d == _T_54[9:0] ? px_buffer_397_g : _GEN_1676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1678 = 10'h18e == _T_54[9:0] ? px_buffer_398_g : _GEN_1677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1679 = 10'h18f == _T_54[9:0] ? px_buffer_399_g : _GEN_1678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1680 = 10'h190 == _T_54[9:0] ? px_buffer_400_g : _GEN_1679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1681 = 10'h191 == _T_54[9:0] ? px_buffer_401_g : _GEN_1680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1682 = 10'h192 == _T_54[9:0] ? px_buffer_402_g : _GEN_1681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1683 = 10'h193 == _T_54[9:0] ? px_buffer_403_g : _GEN_1682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1684 = 10'h194 == _T_54[9:0] ? px_buffer_404_g : _GEN_1683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1685 = 10'h195 == _T_54[9:0] ? px_buffer_405_g : _GEN_1684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1686 = 10'h196 == _T_54[9:0] ? px_buffer_406_g : _GEN_1685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1687 = 10'h197 == _T_54[9:0] ? px_buffer_407_g : _GEN_1686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1688 = 10'h198 == _T_54[9:0] ? px_buffer_408_g : _GEN_1687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1689 = 10'h199 == _T_54[9:0] ? px_buffer_409_g : _GEN_1688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1690 = 10'h19a == _T_54[9:0] ? px_buffer_410_g : _GEN_1689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1691 = 10'h19b == _T_54[9:0] ? px_buffer_411_g : _GEN_1690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1692 = 10'h19c == _T_54[9:0] ? px_buffer_412_g : _GEN_1691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1693 = 10'h19d == _T_54[9:0] ? px_buffer_413_g : _GEN_1692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1694 = 10'h19e == _T_54[9:0] ? px_buffer_414_g : _GEN_1693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1695 = 10'h19f == _T_54[9:0] ? px_buffer_415_g : _GEN_1694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1696 = 10'h1a0 == _T_54[9:0] ? px_buffer_416_g : _GEN_1695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1697 = 10'h1a1 == _T_54[9:0] ? px_buffer_417_g : _GEN_1696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1698 = 10'h1a2 == _T_54[9:0] ? px_buffer_418_g : _GEN_1697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1699 = 10'h1a3 == _T_54[9:0] ? px_buffer_419_g : _GEN_1698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1700 = 10'h1a4 == _T_54[9:0] ? px_buffer_420_g : _GEN_1699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1701 = 10'h1a5 == _T_54[9:0] ? px_buffer_421_g : _GEN_1700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1702 = 10'h1a6 == _T_54[9:0] ? px_buffer_422_g : _GEN_1701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1703 = 10'h1a7 == _T_54[9:0] ? px_buffer_423_g : _GEN_1702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1704 = 10'h1a8 == _T_54[9:0] ? px_buffer_424_g : _GEN_1703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1705 = 10'h1a9 == _T_54[9:0] ? px_buffer_425_g : _GEN_1704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1706 = 10'h1aa == _T_54[9:0] ? px_buffer_426_g : _GEN_1705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1707 = 10'h1ab == _T_54[9:0] ? px_buffer_427_g : _GEN_1706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1708 = 10'h1ac == _T_54[9:0] ? px_buffer_428_g : _GEN_1707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1709 = 10'h1ad == _T_54[9:0] ? px_buffer_429_g : _GEN_1708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1710 = 10'h1ae == _T_54[9:0] ? px_buffer_430_g : _GEN_1709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1711 = 10'h1af == _T_54[9:0] ? px_buffer_431_g : _GEN_1710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1712 = 10'h1b0 == _T_54[9:0] ? px_buffer_432_g : _GEN_1711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1713 = 10'h1b1 == _T_54[9:0] ? px_buffer_433_g : _GEN_1712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1714 = 10'h1b2 == _T_54[9:0] ? px_buffer_434_g : _GEN_1713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1715 = 10'h1b3 == _T_54[9:0] ? px_buffer_435_g : _GEN_1714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1716 = 10'h1b4 == _T_54[9:0] ? px_buffer_436_g : _GEN_1715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1717 = 10'h1b5 == _T_54[9:0] ? px_buffer_437_g : _GEN_1716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1718 = 10'h1b6 == _T_54[9:0] ? px_buffer_438_g : _GEN_1717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1719 = 10'h1b7 == _T_54[9:0] ? px_buffer_439_g : _GEN_1718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1720 = 10'h1b8 == _T_54[9:0] ? px_buffer_440_g : _GEN_1719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1721 = 10'h1b9 == _T_54[9:0] ? px_buffer_441_g : _GEN_1720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1722 = 10'h1ba == _T_54[9:0] ? px_buffer_442_g : _GEN_1721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1723 = 10'h1bb == _T_54[9:0] ? px_buffer_443_g : _GEN_1722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1724 = 10'h1bc == _T_54[9:0] ? px_buffer_444_g : _GEN_1723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1725 = 10'h1bd == _T_54[9:0] ? px_buffer_445_g : _GEN_1724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1726 = 10'h1be == _T_54[9:0] ? px_buffer_446_g : _GEN_1725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1727 = 10'h1bf == _T_54[9:0] ? px_buffer_447_g : _GEN_1726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1728 = 10'h1c0 == _T_54[9:0] ? px_buffer_448_g : _GEN_1727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1729 = 10'h1c1 == _T_54[9:0] ? px_buffer_449_g : _GEN_1728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1730 = 10'h1c2 == _T_54[9:0] ? px_buffer_450_g : _GEN_1729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1731 = 10'h1c3 == _T_54[9:0] ? px_buffer_451_g : _GEN_1730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1732 = 10'h1c4 == _T_54[9:0] ? px_buffer_452_g : _GEN_1731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1733 = 10'h1c5 == _T_54[9:0] ? px_buffer_453_g : _GEN_1732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1734 = 10'h1c6 == _T_54[9:0] ? px_buffer_454_g : _GEN_1733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1735 = 10'h1c7 == _T_54[9:0] ? px_buffer_455_g : _GEN_1734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1736 = 10'h1c8 == _T_54[9:0] ? px_buffer_456_g : _GEN_1735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1737 = 10'h1c9 == _T_54[9:0] ? px_buffer_457_g : _GEN_1736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1738 = 10'h1ca == _T_54[9:0] ? px_buffer_458_g : _GEN_1737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1739 = 10'h1cb == _T_54[9:0] ? px_buffer_459_g : _GEN_1738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1740 = 10'h1cc == _T_54[9:0] ? px_buffer_460_g : _GEN_1739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1741 = 10'h1cd == _T_54[9:0] ? px_buffer_461_g : _GEN_1740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1742 = 10'h1ce == _T_54[9:0] ? px_buffer_462_g : _GEN_1741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1743 = 10'h1cf == _T_54[9:0] ? px_buffer_463_g : _GEN_1742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1744 = 10'h1d0 == _T_54[9:0] ? px_buffer_464_g : _GEN_1743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1745 = 10'h1d1 == _T_54[9:0] ? px_buffer_465_g : _GEN_1744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1746 = 10'h1d2 == _T_54[9:0] ? px_buffer_466_g : _GEN_1745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1747 = 10'h1d3 == _T_54[9:0] ? px_buffer_467_g : _GEN_1746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1748 = 10'h1d4 == _T_54[9:0] ? px_buffer_468_g : _GEN_1747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1749 = 10'h1d5 == _T_54[9:0] ? px_buffer_469_g : _GEN_1748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1750 = 10'h1d6 == _T_54[9:0] ? px_buffer_470_g : _GEN_1749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1751 = 10'h1d7 == _T_54[9:0] ? px_buffer_471_g : _GEN_1750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1752 = 10'h1d8 == _T_54[9:0] ? px_buffer_472_g : _GEN_1751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1753 = 10'h1d9 == _T_54[9:0] ? px_buffer_473_g : _GEN_1752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1754 = 10'h1da == _T_54[9:0] ? px_buffer_474_g : _GEN_1753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1755 = 10'h1db == _T_54[9:0] ? px_buffer_475_g : _GEN_1754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1756 = 10'h1dc == _T_54[9:0] ? px_buffer_476_g : _GEN_1755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1757 = 10'h1dd == _T_54[9:0] ? px_buffer_477_g : _GEN_1756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1758 = 10'h1de == _T_54[9:0] ? px_buffer_478_g : _GEN_1757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1759 = 10'h1df == _T_54[9:0] ? px_buffer_479_g : _GEN_1758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1760 = 10'h1e0 == _T_54[9:0] ? px_buffer_480_g : _GEN_1759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1761 = 10'h1e1 == _T_54[9:0] ? px_buffer_481_g : _GEN_1760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1762 = 10'h1e2 == _T_54[9:0] ? px_buffer_482_g : _GEN_1761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1763 = 10'h1e3 == _T_54[9:0] ? px_buffer_483_g : _GEN_1762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1764 = 10'h1e4 == _T_54[9:0] ? px_buffer_484_g : _GEN_1763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1765 = 10'h1e5 == _T_54[9:0] ? px_buffer_485_g : _GEN_1764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1766 = 10'h1e6 == _T_54[9:0] ? px_buffer_486_g : _GEN_1765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1767 = 10'h1e7 == _T_54[9:0] ? px_buffer_487_g : _GEN_1766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1768 = 10'h1e8 == _T_54[9:0] ? px_buffer_488_g : _GEN_1767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1769 = 10'h1e9 == _T_54[9:0] ? px_buffer_489_g : _GEN_1768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1770 = 10'h1ea == _T_54[9:0] ? px_buffer_490_g : _GEN_1769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1771 = 10'h1eb == _T_54[9:0] ? px_buffer_491_g : _GEN_1770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1772 = 10'h1ec == _T_54[9:0] ? px_buffer_492_g : _GEN_1771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1773 = 10'h1ed == _T_54[9:0] ? px_buffer_493_g : _GEN_1772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1774 = 10'h1ee == _T_54[9:0] ? px_buffer_494_g : _GEN_1773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1775 = 10'h1ef == _T_54[9:0] ? px_buffer_495_g : _GEN_1774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1776 = 10'h1f0 == _T_54[9:0] ? px_buffer_496_g : _GEN_1775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1777 = 10'h1f1 == _T_54[9:0] ? px_buffer_497_g : _GEN_1776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1778 = 10'h1f2 == _T_54[9:0] ? px_buffer_498_g : _GEN_1777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1779 = 10'h1f3 == _T_54[9:0] ? px_buffer_499_g : _GEN_1778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1780 = 10'h1f4 == _T_54[9:0] ? px_buffer_500_g : _GEN_1779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1781 = 10'h1f5 == _T_54[9:0] ? px_buffer_501_g : _GEN_1780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1782 = 10'h1f6 == _T_54[9:0] ? px_buffer_502_g : _GEN_1781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1783 = 10'h1f7 == _T_54[9:0] ? px_buffer_503_g : _GEN_1782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1784 = 10'h1f8 == _T_54[9:0] ? px_buffer_504_g : _GEN_1783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1785 = 10'h1f9 == _T_54[9:0] ? px_buffer_505_g : _GEN_1784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1786 = 10'h1fa == _T_54[9:0] ? px_buffer_506_g : _GEN_1785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1787 = 10'h1fb == _T_54[9:0] ? px_buffer_507_g : _GEN_1786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1788 = 10'h1fc == _T_54[9:0] ? px_buffer_508_g : _GEN_1787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1789 = 10'h1fd == _T_54[9:0] ? px_buffer_509_g : _GEN_1788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1790 = 10'h1fe == _T_54[9:0] ? px_buffer_510_g : _GEN_1789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1791 = 10'h1ff == _T_54[9:0] ? px_buffer_511_g : _GEN_1790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1792 = 10'h200 == _T_54[9:0] ? px_buffer_512_g : _GEN_1791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1793 = 10'h201 == _T_54[9:0] ? px_buffer_513_g : _GEN_1792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1794 = 10'h202 == _T_54[9:0] ? px_buffer_514_g : _GEN_1793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1795 = 10'h203 == _T_54[9:0] ? px_buffer_515_g : _GEN_1794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1796 = 10'h204 == _T_54[9:0] ? px_buffer_516_g : _GEN_1795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1797 = 10'h205 == _T_54[9:0] ? px_buffer_517_g : _GEN_1796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1798 = 10'h206 == _T_54[9:0] ? px_buffer_518_g : _GEN_1797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1799 = 10'h207 == _T_54[9:0] ? px_buffer_519_g : _GEN_1798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1800 = 10'h208 == _T_54[9:0] ? px_buffer_520_g : _GEN_1799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1801 = 10'h209 == _T_54[9:0] ? px_buffer_521_g : _GEN_1800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1802 = 10'h20a == _T_54[9:0] ? px_buffer_522_g : _GEN_1801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1803 = 10'h20b == _T_54[9:0] ? px_buffer_523_g : _GEN_1802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1804 = 10'h20c == _T_54[9:0] ? px_buffer_524_g : _GEN_1803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1805 = 10'h20d == _T_54[9:0] ? px_buffer_525_g : _GEN_1804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1806 = 10'h20e == _T_54[9:0] ? px_buffer_526_g : _GEN_1805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1807 = 10'h20f == _T_54[9:0] ? px_buffer_527_g : _GEN_1806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1808 = 10'h210 == _T_54[9:0] ? px_buffer_528_g : _GEN_1807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1809 = 10'h211 == _T_54[9:0] ? px_buffer_529_g : _GEN_1808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1810 = 10'h212 == _T_54[9:0] ? px_buffer_530_g : _GEN_1809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1811 = 10'h213 == _T_54[9:0] ? px_buffer_531_g : _GEN_1810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1812 = 10'h214 == _T_54[9:0] ? px_buffer_532_g : _GEN_1811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1813 = 10'h215 == _T_54[9:0] ? px_buffer_533_g : _GEN_1812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1814 = 10'h216 == _T_54[9:0] ? px_buffer_534_g : _GEN_1813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1815 = 10'h217 == _T_54[9:0] ? px_buffer_535_g : _GEN_1814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1816 = 10'h218 == _T_54[9:0] ? px_buffer_536_g : _GEN_1815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1817 = 10'h219 == _T_54[9:0] ? px_buffer_537_g : _GEN_1816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1818 = 10'h21a == _T_54[9:0] ? px_buffer_538_g : _GEN_1817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1819 = 10'h21b == _T_54[9:0] ? px_buffer_539_g : _GEN_1818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1820 = 10'h21c == _T_54[9:0] ? px_buffer_540_g : _GEN_1819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1821 = 10'h21d == _T_54[9:0] ? px_buffer_541_g : _GEN_1820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1822 = 10'h21e == _T_54[9:0] ? px_buffer_542_g : _GEN_1821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1823 = 10'h21f == _T_54[9:0] ? px_buffer_543_g : _GEN_1822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1824 = 10'h220 == _T_54[9:0] ? px_buffer_544_g : _GEN_1823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1825 = 10'h221 == _T_54[9:0] ? px_buffer_545_g : _GEN_1824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1826 = 10'h222 == _T_54[9:0] ? px_buffer_546_g : _GEN_1825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1827 = 10'h223 == _T_54[9:0] ? px_buffer_547_g : _GEN_1826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1828 = 10'h224 == _T_54[9:0] ? px_buffer_548_g : _GEN_1827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1829 = 10'h225 == _T_54[9:0] ? px_buffer_549_g : _GEN_1828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1830 = 10'h226 == _T_54[9:0] ? px_buffer_550_g : _GEN_1829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1831 = 10'h227 == _T_54[9:0] ? px_buffer_551_g : _GEN_1830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1832 = 10'h228 == _T_54[9:0] ? px_buffer_552_g : _GEN_1831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1833 = 10'h229 == _T_54[9:0] ? px_buffer_553_g : _GEN_1832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1834 = 10'h22a == _T_54[9:0] ? px_buffer_554_g : _GEN_1833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1835 = 10'h22b == _T_54[9:0] ? px_buffer_555_g : _GEN_1834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1836 = 10'h22c == _T_54[9:0] ? px_buffer_556_g : _GEN_1835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1837 = 10'h22d == _T_54[9:0] ? px_buffer_557_g : _GEN_1836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1838 = 10'h22e == _T_54[9:0] ? px_buffer_558_g : _GEN_1837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1839 = 10'h22f == _T_54[9:0] ? px_buffer_559_g : _GEN_1838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1840 = 10'h230 == _T_54[9:0] ? px_buffer_560_g : _GEN_1839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1841 = 10'h231 == _T_54[9:0] ? px_buffer_561_g : _GEN_1840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1842 = 10'h232 == _T_54[9:0] ? px_buffer_562_g : _GEN_1841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1843 = 10'h233 == _T_54[9:0] ? px_buffer_563_g : _GEN_1842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1844 = 10'h234 == _T_54[9:0] ? px_buffer_564_g : _GEN_1843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1845 = 10'h235 == _T_54[9:0] ? px_buffer_565_g : _GEN_1844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1846 = 10'h236 == _T_54[9:0] ? px_buffer_566_g : _GEN_1845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1847 = 10'h237 == _T_54[9:0] ? px_buffer_567_g : _GEN_1846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1848 = 10'h238 == _T_54[9:0] ? px_buffer_568_g : _GEN_1847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1849 = 10'h239 == _T_54[9:0] ? px_buffer_569_g : _GEN_1848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1850 = 10'h23a == _T_54[9:0] ? px_buffer_570_g : _GEN_1849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1851 = 10'h23b == _T_54[9:0] ? px_buffer_571_g : _GEN_1850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1852 = 10'h23c == _T_54[9:0] ? px_buffer_572_g : _GEN_1851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1853 = 10'h23d == _T_54[9:0] ? px_buffer_573_g : _GEN_1852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1854 = 10'h23e == _T_54[9:0] ? px_buffer_574_g : _GEN_1853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1855 = 10'h23f == _T_54[9:0] ? px_buffer_575_g : _GEN_1854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1856 = 10'h240 == _T_54[9:0] ? px_buffer_576_g : _GEN_1855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1857 = 10'h241 == _T_54[9:0] ? px_buffer_577_g : _GEN_1856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1858 = 10'h242 == _T_54[9:0] ? px_buffer_578_g : _GEN_1857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1859 = 10'h243 == _T_54[9:0] ? px_buffer_579_g : _GEN_1858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1860 = 10'h244 == _T_54[9:0] ? px_buffer_580_g : _GEN_1859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1861 = 10'h245 == _T_54[9:0] ? px_buffer_581_g : _GEN_1860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1862 = 10'h246 == _T_54[9:0] ? px_buffer_582_g : _GEN_1861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1863 = 10'h247 == _T_54[9:0] ? px_buffer_583_g : _GEN_1862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1864 = 10'h248 == _T_54[9:0] ? px_buffer_584_g : _GEN_1863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1865 = 10'h249 == _T_54[9:0] ? px_buffer_585_g : _GEN_1864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1866 = 10'h24a == _T_54[9:0] ? px_buffer_586_g : _GEN_1865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1867 = 10'h24b == _T_54[9:0] ? px_buffer_587_g : _GEN_1866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1868 = 10'h24c == _T_54[9:0] ? px_buffer_588_g : _GEN_1867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1869 = 10'h24d == _T_54[9:0] ? px_buffer_589_g : _GEN_1868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1870 = 10'h24e == _T_54[9:0] ? px_buffer_590_g : _GEN_1869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1871 = 10'h24f == _T_54[9:0] ? px_buffer_591_g : _GEN_1870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1872 = 10'h250 == _T_54[9:0] ? px_buffer_592_g : _GEN_1871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1873 = 10'h251 == _T_54[9:0] ? px_buffer_593_g : _GEN_1872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1874 = 10'h252 == _T_54[9:0] ? px_buffer_594_g : _GEN_1873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1875 = 10'h253 == _T_54[9:0] ? px_buffer_595_g : _GEN_1874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1876 = 10'h254 == _T_54[9:0] ? px_buffer_596_g : _GEN_1875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1877 = 10'h255 == _T_54[9:0] ? px_buffer_597_g : _GEN_1876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1878 = 10'h256 == _T_54[9:0] ? px_buffer_598_g : _GEN_1877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1879 = 10'h257 == _T_54[9:0] ? px_buffer_599_g : _GEN_1878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1880 = 10'h258 == _T_54[9:0] ? px_buffer_600_g : _GEN_1879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1881 = 10'h259 == _T_54[9:0] ? px_buffer_601_g : _GEN_1880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1882 = 10'h25a == _T_54[9:0] ? px_buffer_602_g : _GEN_1881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1883 = 10'h25b == _T_54[9:0] ? px_buffer_603_g : _GEN_1882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1884 = 10'h25c == _T_54[9:0] ? px_buffer_604_g : _GEN_1883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1885 = 10'h25d == _T_54[9:0] ? px_buffer_605_g : _GEN_1884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1886 = 10'h25e == _T_54[9:0] ? px_buffer_606_g : _GEN_1885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1887 = 10'h25f == _T_54[9:0] ? px_buffer_607_g : _GEN_1886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1888 = 10'h260 == _T_54[9:0] ? px_buffer_608_g : _GEN_1887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1889 = 10'h261 == _T_54[9:0] ? px_buffer_609_g : _GEN_1888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1890 = 10'h262 == _T_54[9:0] ? px_buffer_610_g : _GEN_1889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1891 = 10'h263 == _T_54[9:0] ? px_buffer_611_g : _GEN_1890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1892 = 10'h264 == _T_54[9:0] ? px_buffer_612_g : _GEN_1891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1893 = 10'h265 == _T_54[9:0] ? px_buffer_613_g : _GEN_1892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1894 = 10'h266 == _T_54[9:0] ? px_buffer_614_g : _GEN_1893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1895 = 10'h267 == _T_54[9:0] ? px_buffer_615_g : _GEN_1894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1896 = 10'h268 == _T_54[9:0] ? px_buffer_616_g : _GEN_1895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1897 = 10'h269 == _T_54[9:0] ? px_buffer_617_g : _GEN_1896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1898 = 10'h26a == _T_54[9:0] ? px_buffer_618_g : _GEN_1897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1899 = 10'h26b == _T_54[9:0] ? px_buffer_619_g : _GEN_1898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1900 = 10'h26c == _T_54[9:0] ? px_buffer_620_g : _GEN_1899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1901 = 10'h26d == _T_54[9:0] ? px_buffer_621_g : _GEN_1900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1902 = 10'h26e == _T_54[9:0] ? px_buffer_622_g : _GEN_1901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1903 = 10'h26f == _T_54[9:0] ? px_buffer_623_g : _GEN_1902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1904 = 10'h270 == _T_54[9:0] ? px_buffer_624_g : _GEN_1903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1905 = 10'h271 == _T_54[9:0] ? px_buffer_625_g : _GEN_1904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1906 = 10'h272 == _T_54[9:0] ? px_buffer_626_g : _GEN_1905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1907 = 10'h273 == _T_54[9:0] ? px_buffer_627_g : _GEN_1906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1908 = 10'h274 == _T_54[9:0] ? px_buffer_628_g : _GEN_1907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1909 = 10'h275 == _T_54[9:0] ? px_buffer_629_g : _GEN_1908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1910 = 10'h276 == _T_54[9:0] ? px_buffer_630_g : _GEN_1909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1911 = 10'h277 == _T_54[9:0] ? px_buffer_631_g : _GEN_1910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1912 = 10'h278 == _T_54[9:0] ? px_buffer_632_g : _GEN_1911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1913 = 10'h279 == _T_54[9:0] ? px_buffer_633_g : _GEN_1912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1914 = 10'h27a == _T_54[9:0] ? px_buffer_634_g : _GEN_1913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1915 = 10'h27b == _T_54[9:0] ? px_buffer_635_g : _GEN_1914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1916 = 10'h27c == _T_54[9:0] ? px_buffer_636_g : _GEN_1915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1917 = 10'h27d == _T_54[9:0] ? px_buffer_637_g : _GEN_1916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1918 = 10'h27e == _T_54[9:0] ? px_buffer_638_g : _GEN_1917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1919 = 10'h27f == _T_54[9:0] ? px_buffer_639_g : _GEN_1918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _T_75 = {1'h0,_GEN_1919}; // @[EdgeDetect.scala 56:51]
  wire [8:0] _T_77 = {1'h0,io_px_in_g}; // @[EdgeDetect.scala 56:81]
  wire [8:0] _T_80 = $signed(_T_75) - $signed(_T_77); // @[EdgeDetect.scala 56:58]
  wire [7:0] _GEN_1921 = 10'h1 == io_x[9:0] ? px_buffer_1_g : px_buffer_0_g; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1922 = 10'h2 == io_x[9:0] ? px_buffer_2_g : _GEN_1921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1923 = 10'h3 == io_x[9:0] ? px_buffer_3_g : _GEN_1922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1924 = 10'h4 == io_x[9:0] ? px_buffer_4_g : _GEN_1923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1925 = 10'h5 == io_x[9:0] ? px_buffer_5_g : _GEN_1924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1926 = 10'h6 == io_x[9:0] ? px_buffer_6_g : _GEN_1925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1927 = 10'h7 == io_x[9:0] ? px_buffer_7_g : _GEN_1926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1928 = 10'h8 == io_x[9:0] ? px_buffer_8_g : _GEN_1927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1929 = 10'h9 == io_x[9:0] ? px_buffer_9_g : _GEN_1928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1930 = 10'ha == io_x[9:0] ? px_buffer_10_g : _GEN_1929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1931 = 10'hb == io_x[9:0] ? px_buffer_11_g : _GEN_1930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1932 = 10'hc == io_x[9:0] ? px_buffer_12_g : _GEN_1931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1933 = 10'hd == io_x[9:0] ? px_buffer_13_g : _GEN_1932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1934 = 10'he == io_x[9:0] ? px_buffer_14_g : _GEN_1933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1935 = 10'hf == io_x[9:0] ? px_buffer_15_g : _GEN_1934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1936 = 10'h10 == io_x[9:0] ? px_buffer_16_g : _GEN_1935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1937 = 10'h11 == io_x[9:0] ? px_buffer_17_g : _GEN_1936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1938 = 10'h12 == io_x[9:0] ? px_buffer_18_g : _GEN_1937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1939 = 10'h13 == io_x[9:0] ? px_buffer_19_g : _GEN_1938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1940 = 10'h14 == io_x[9:0] ? px_buffer_20_g : _GEN_1939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1941 = 10'h15 == io_x[9:0] ? px_buffer_21_g : _GEN_1940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1942 = 10'h16 == io_x[9:0] ? px_buffer_22_g : _GEN_1941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1943 = 10'h17 == io_x[9:0] ? px_buffer_23_g : _GEN_1942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1944 = 10'h18 == io_x[9:0] ? px_buffer_24_g : _GEN_1943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1945 = 10'h19 == io_x[9:0] ? px_buffer_25_g : _GEN_1944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1946 = 10'h1a == io_x[9:0] ? px_buffer_26_g : _GEN_1945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1947 = 10'h1b == io_x[9:0] ? px_buffer_27_g : _GEN_1946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1948 = 10'h1c == io_x[9:0] ? px_buffer_28_g : _GEN_1947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1949 = 10'h1d == io_x[9:0] ? px_buffer_29_g : _GEN_1948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1950 = 10'h1e == io_x[9:0] ? px_buffer_30_g : _GEN_1949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1951 = 10'h1f == io_x[9:0] ? px_buffer_31_g : _GEN_1950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1952 = 10'h20 == io_x[9:0] ? px_buffer_32_g : _GEN_1951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1953 = 10'h21 == io_x[9:0] ? px_buffer_33_g : _GEN_1952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1954 = 10'h22 == io_x[9:0] ? px_buffer_34_g : _GEN_1953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1955 = 10'h23 == io_x[9:0] ? px_buffer_35_g : _GEN_1954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1956 = 10'h24 == io_x[9:0] ? px_buffer_36_g : _GEN_1955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1957 = 10'h25 == io_x[9:0] ? px_buffer_37_g : _GEN_1956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1958 = 10'h26 == io_x[9:0] ? px_buffer_38_g : _GEN_1957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1959 = 10'h27 == io_x[9:0] ? px_buffer_39_g : _GEN_1958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1960 = 10'h28 == io_x[9:0] ? px_buffer_40_g : _GEN_1959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1961 = 10'h29 == io_x[9:0] ? px_buffer_41_g : _GEN_1960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1962 = 10'h2a == io_x[9:0] ? px_buffer_42_g : _GEN_1961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1963 = 10'h2b == io_x[9:0] ? px_buffer_43_g : _GEN_1962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1964 = 10'h2c == io_x[9:0] ? px_buffer_44_g : _GEN_1963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1965 = 10'h2d == io_x[9:0] ? px_buffer_45_g : _GEN_1964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1966 = 10'h2e == io_x[9:0] ? px_buffer_46_g : _GEN_1965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1967 = 10'h2f == io_x[9:0] ? px_buffer_47_g : _GEN_1966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1968 = 10'h30 == io_x[9:0] ? px_buffer_48_g : _GEN_1967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1969 = 10'h31 == io_x[9:0] ? px_buffer_49_g : _GEN_1968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1970 = 10'h32 == io_x[9:0] ? px_buffer_50_g : _GEN_1969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1971 = 10'h33 == io_x[9:0] ? px_buffer_51_g : _GEN_1970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1972 = 10'h34 == io_x[9:0] ? px_buffer_52_g : _GEN_1971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1973 = 10'h35 == io_x[9:0] ? px_buffer_53_g : _GEN_1972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1974 = 10'h36 == io_x[9:0] ? px_buffer_54_g : _GEN_1973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1975 = 10'h37 == io_x[9:0] ? px_buffer_55_g : _GEN_1974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1976 = 10'h38 == io_x[9:0] ? px_buffer_56_g : _GEN_1975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1977 = 10'h39 == io_x[9:0] ? px_buffer_57_g : _GEN_1976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1978 = 10'h3a == io_x[9:0] ? px_buffer_58_g : _GEN_1977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1979 = 10'h3b == io_x[9:0] ? px_buffer_59_g : _GEN_1978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1980 = 10'h3c == io_x[9:0] ? px_buffer_60_g : _GEN_1979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1981 = 10'h3d == io_x[9:0] ? px_buffer_61_g : _GEN_1980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1982 = 10'h3e == io_x[9:0] ? px_buffer_62_g : _GEN_1981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1983 = 10'h3f == io_x[9:0] ? px_buffer_63_g : _GEN_1982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1984 = 10'h40 == io_x[9:0] ? px_buffer_64_g : _GEN_1983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1985 = 10'h41 == io_x[9:0] ? px_buffer_65_g : _GEN_1984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1986 = 10'h42 == io_x[9:0] ? px_buffer_66_g : _GEN_1985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1987 = 10'h43 == io_x[9:0] ? px_buffer_67_g : _GEN_1986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1988 = 10'h44 == io_x[9:0] ? px_buffer_68_g : _GEN_1987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1989 = 10'h45 == io_x[9:0] ? px_buffer_69_g : _GEN_1988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1990 = 10'h46 == io_x[9:0] ? px_buffer_70_g : _GEN_1989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1991 = 10'h47 == io_x[9:0] ? px_buffer_71_g : _GEN_1990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1992 = 10'h48 == io_x[9:0] ? px_buffer_72_g : _GEN_1991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1993 = 10'h49 == io_x[9:0] ? px_buffer_73_g : _GEN_1992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1994 = 10'h4a == io_x[9:0] ? px_buffer_74_g : _GEN_1993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1995 = 10'h4b == io_x[9:0] ? px_buffer_75_g : _GEN_1994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1996 = 10'h4c == io_x[9:0] ? px_buffer_76_g : _GEN_1995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1997 = 10'h4d == io_x[9:0] ? px_buffer_77_g : _GEN_1996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1998 = 10'h4e == io_x[9:0] ? px_buffer_78_g : _GEN_1997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1999 = 10'h4f == io_x[9:0] ? px_buffer_79_g : _GEN_1998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2000 = 10'h50 == io_x[9:0] ? px_buffer_80_g : _GEN_1999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2001 = 10'h51 == io_x[9:0] ? px_buffer_81_g : _GEN_2000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2002 = 10'h52 == io_x[9:0] ? px_buffer_82_g : _GEN_2001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2003 = 10'h53 == io_x[9:0] ? px_buffer_83_g : _GEN_2002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2004 = 10'h54 == io_x[9:0] ? px_buffer_84_g : _GEN_2003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2005 = 10'h55 == io_x[9:0] ? px_buffer_85_g : _GEN_2004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2006 = 10'h56 == io_x[9:0] ? px_buffer_86_g : _GEN_2005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2007 = 10'h57 == io_x[9:0] ? px_buffer_87_g : _GEN_2006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2008 = 10'h58 == io_x[9:0] ? px_buffer_88_g : _GEN_2007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2009 = 10'h59 == io_x[9:0] ? px_buffer_89_g : _GEN_2008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2010 = 10'h5a == io_x[9:0] ? px_buffer_90_g : _GEN_2009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2011 = 10'h5b == io_x[9:0] ? px_buffer_91_g : _GEN_2010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2012 = 10'h5c == io_x[9:0] ? px_buffer_92_g : _GEN_2011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2013 = 10'h5d == io_x[9:0] ? px_buffer_93_g : _GEN_2012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2014 = 10'h5e == io_x[9:0] ? px_buffer_94_g : _GEN_2013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2015 = 10'h5f == io_x[9:0] ? px_buffer_95_g : _GEN_2014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2016 = 10'h60 == io_x[9:0] ? px_buffer_96_g : _GEN_2015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2017 = 10'h61 == io_x[9:0] ? px_buffer_97_g : _GEN_2016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2018 = 10'h62 == io_x[9:0] ? px_buffer_98_g : _GEN_2017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2019 = 10'h63 == io_x[9:0] ? px_buffer_99_g : _GEN_2018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2020 = 10'h64 == io_x[9:0] ? px_buffer_100_g : _GEN_2019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2021 = 10'h65 == io_x[9:0] ? px_buffer_101_g : _GEN_2020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2022 = 10'h66 == io_x[9:0] ? px_buffer_102_g : _GEN_2021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2023 = 10'h67 == io_x[9:0] ? px_buffer_103_g : _GEN_2022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2024 = 10'h68 == io_x[9:0] ? px_buffer_104_g : _GEN_2023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2025 = 10'h69 == io_x[9:0] ? px_buffer_105_g : _GEN_2024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2026 = 10'h6a == io_x[9:0] ? px_buffer_106_g : _GEN_2025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2027 = 10'h6b == io_x[9:0] ? px_buffer_107_g : _GEN_2026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2028 = 10'h6c == io_x[9:0] ? px_buffer_108_g : _GEN_2027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2029 = 10'h6d == io_x[9:0] ? px_buffer_109_g : _GEN_2028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2030 = 10'h6e == io_x[9:0] ? px_buffer_110_g : _GEN_2029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2031 = 10'h6f == io_x[9:0] ? px_buffer_111_g : _GEN_2030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2032 = 10'h70 == io_x[9:0] ? px_buffer_112_g : _GEN_2031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2033 = 10'h71 == io_x[9:0] ? px_buffer_113_g : _GEN_2032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2034 = 10'h72 == io_x[9:0] ? px_buffer_114_g : _GEN_2033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2035 = 10'h73 == io_x[9:0] ? px_buffer_115_g : _GEN_2034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2036 = 10'h74 == io_x[9:0] ? px_buffer_116_g : _GEN_2035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2037 = 10'h75 == io_x[9:0] ? px_buffer_117_g : _GEN_2036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2038 = 10'h76 == io_x[9:0] ? px_buffer_118_g : _GEN_2037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2039 = 10'h77 == io_x[9:0] ? px_buffer_119_g : _GEN_2038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2040 = 10'h78 == io_x[9:0] ? px_buffer_120_g : _GEN_2039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2041 = 10'h79 == io_x[9:0] ? px_buffer_121_g : _GEN_2040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2042 = 10'h7a == io_x[9:0] ? px_buffer_122_g : _GEN_2041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2043 = 10'h7b == io_x[9:0] ? px_buffer_123_g : _GEN_2042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2044 = 10'h7c == io_x[9:0] ? px_buffer_124_g : _GEN_2043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2045 = 10'h7d == io_x[9:0] ? px_buffer_125_g : _GEN_2044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2046 = 10'h7e == io_x[9:0] ? px_buffer_126_g : _GEN_2045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2047 = 10'h7f == io_x[9:0] ? px_buffer_127_g : _GEN_2046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2048 = 10'h80 == io_x[9:0] ? px_buffer_128_g : _GEN_2047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2049 = 10'h81 == io_x[9:0] ? px_buffer_129_g : _GEN_2048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2050 = 10'h82 == io_x[9:0] ? px_buffer_130_g : _GEN_2049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2051 = 10'h83 == io_x[9:0] ? px_buffer_131_g : _GEN_2050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2052 = 10'h84 == io_x[9:0] ? px_buffer_132_g : _GEN_2051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2053 = 10'h85 == io_x[9:0] ? px_buffer_133_g : _GEN_2052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2054 = 10'h86 == io_x[9:0] ? px_buffer_134_g : _GEN_2053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2055 = 10'h87 == io_x[9:0] ? px_buffer_135_g : _GEN_2054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2056 = 10'h88 == io_x[9:0] ? px_buffer_136_g : _GEN_2055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2057 = 10'h89 == io_x[9:0] ? px_buffer_137_g : _GEN_2056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2058 = 10'h8a == io_x[9:0] ? px_buffer_138_g : _GEN_2057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2059 = 10'h8b == io_x[9:0] ? px_buffer_139_g : _GEN_2058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2060 = 10'h8c == io_x[9:0] ? px_buffer_140_g : _GEN_2059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2061 = 10'h8d == io_x[9:0] ? px_buffer_141_g : _GEN_2060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2062 = 10'h8e == io_x[9:0] ? px_buffer_142_g : _GEN_2061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2063 = 10'h8f == io_x[9:0] ? px_buffer_143_g : _GEN_2062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2064 = 10'h90 == io_x[9:0] ? px_buffer_144_g : _GEN_2063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2065 = 10'h91 == io_x[9:0] ? px_buffer_145_g : _GEN_2064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2066 = 10'h92 == io_x[9:0] ? px_buffer_146_g : _GEN_2065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2067 = 10'h93 == io_x[9:0] ? px_buffer_147_g : _GEN_2066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2068 = 10'h94 == io_x[9:0] ? px_buffer_148_g : _GEN_2067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2069 = 10'h95 == io_x[9:0] ? px_buffer_149_g : _GEN_2068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2070 = 10'h96 == io_x[9:0] ? px_buffer_150_g : _GEN_2069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2071 = 10'h97 == io_x[9:0] ? px_buffer_151_g : _GEN_2070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2072 = 10'h98 == io_x[9:0] ? px_buffer_152_g : _GEN_2071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2073 = 10'h99 == io_x[9:0] ? px_buffer_153_g : _GEN_2072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2074 = 10'h9a == io_x[9:0] ? px_buffer_154_g : _GEN_2073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2075 = 10'h9b == io_x[9:0] ? px_buffer_155_g : _GEN_2074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2076 = 10'h9c == io_x[9:0] ? px_buffer_156_g : _GEN_2075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2077 = 10'h9d == io_x[9:0] ? px_buffer_157_g : _GEN_2076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2078 = 10'h9e == io_x[9:0] ? px_buffer_158_g : _GEN_2077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2079 = 10'h9f == io_x[9:0] ? px_buffer_159_g : _GEN_2078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2080 = 10'ha0 == io_x[9:0] ? px_buffer_160_g : _GEN_2079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2081 = 10'ha1 == io_x[9:0] ? px_buffer_161_g : _GEN_2080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2082 = 10'ha2 == io_x[9:0] ? px_buffer_162_g : _GEN_2081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2083 = 10'ha3 == io_x[9:0] ? px_buffer_163_g : _GEN_2082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2084 = 10'ha4 == io_x[9:0] ? px_buffer_164_g : _GEN_2083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2085 = 10'ha5 == io_x[9:0] ? px_buffer_165_g : _GEN_2084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2086 = 10'ha6 == io_x[9:0] ? px_buffer_166_g : _GEN_2085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2087 = 10'ha7 == io_x[9:0] ? px_buffer_167_g : _GEN_2086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2088 = 10'ha8 == io_x[9:0] ? px_buffer_168_g : _GEN_2087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2089 = 10'ha9 == io_x[9:0] ? px_buffer_169_g : _GEN_2088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2090 = 10'haa == io_x[9:0] ? px_buffer_170_g : _GEN_2089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2091 = 10'hab == io_x[9:0] ? px_buffer_171_g : _GEN_2090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2092 = 10'hac == io_x[9:0] ? px_buffer_172_g : _GEN_2091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2093 = 10'had == io_x[9:0] ? px_buffer_173_g : _GEN_2092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2094 = 10'hae == io_x[9:0] ? px_buffer_174_g : _GEN_2093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2095 = 10'haf == io_x[9:0] ? px_buffer_175_g : _GEN_2094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2096 = 10'hb0 == io_x[9:0] ? px_buffer_176_g : _GEN_2095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2097 = 10'hb1 == io_x[9:0] ? px_buffer_177_g : _GEN_2096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2098 = 10'hb2 == io_x[9:0] ? px_buffer_178_g : _GEN_2097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2099 = 10'hb3 == io_x[9:0] ? px_buffer_179_g : _GEN_2098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2100 = 10'hb4 == io_x[9:0] ? px_buffer_180_g : _GEN_2099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2101 = 10'hb5 == io_x[9:0] ? px_buffer_181_g : _GEN_2100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2102 = 10'hb6 == io_x[9:0] ? px_buffer_182_g : _GEN_2101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2103 = 10'hb7 == io_x[9:0] ? px_buffer_183_g : _GEN_2102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2104 = 10'hb8 == io_x[9:0] ? px_buffer_184_g : _GEN_2103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2105 = 10'hb9 == io_x[9:0] ? px_buffer_185_g : _GEN_2104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2106 = 10'hba == io_x[9:0] ? px_buffer_186_g : _GEN_2105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2107 = 10'hbb == io_x[9:0] ? px_buffer_187_g : _GEN_2106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2108 = 10'hbc == io_x[9:0] ? px_buffer_188_g : _GEN_2107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2109 = 10'hbd == io_x[9:0] ? px_buffer_189_g : _GEN_2108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2110 = 10'hbe == io_x[9:0] ? px_buffer_190_g : _GEN_2109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2111 = 10'hbf == io_x[9:0] ? px_buffer_191_g : _GEN_2110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2112 = 10'hc0 == io_x[9:0] ? px_buffer_192_g : _GEN_2111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2113 = 10'hc1 == io_x[9:0] ? px_buffer_193_g : _GEN_2112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2114 = 10'hc2 == io_x[9:0] ? px_buffer_194_g : _GEN_2113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2115 = 10'hc3 == io_x[9:0] ? px_buffer_195_g : _GEN_2114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2116 = 10'hc4 == io_x[9:0] ? px_buffer_196_g : _GEN_2115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2117 = 10'hc5 == io_x[9:0] ? px_buffer_197_g : _GEN_2116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2118 = 10'hc6 == io_x[9:0] ? px_buffer_198_g : _GEN_2117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2119 = 10'hc7 == io_x[9:0] ? px_buffer_199_g : _GEN_2118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2120 = 10'hc8 == io_x[9:0] ? px_buffer_200_g : _GEN_2119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2121 = 10'hc9 == io_x[9:0] ? px_buffer_201_g : _GEN_2120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2122 = 10'hca == io_x[9:0] ? px_buffer_202_g : _GEN_2121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2123 = 10'hcb == io_x[9:0] ? px_buffer_203_g : _GEN_2122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2124 = 10'hcc == io_x[9:0] ? px_buffer_204_g : _GEN_2123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2125 = 10'hcd == io_x[9:0] ? px_buffer_205_g : _GEN_2124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2126 = 10'hce == io_x[9:0] ? px_buffer_206_g : _GEN_2125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2127 = 10'hcf == io_x[9:0] ? px_buffer_207_g : _GEN_2126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2128 = 10'hd0 == io_x[9:0] ? px_buffer_208_g : _GEN_2127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2129 = 10'hd1 == io_x[9:0] ? px_buffer_209_g : _GEN_2128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2130 = 10'hd2 == io_x[9:0] ? px_buffer_210_g : _GEN_2129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2131 = 10'hd3 == io_x[9:0] ? px_buffer_211_g : _GEN_2130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2132 = 10'hd4 == io_x[9:0] ? px_buffer_212_g : _GEN_2131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2133 = 10'hd5 == io_x[9:0] ? px_buffer_213_g : _GEN_2132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2134 = 10'hd6 == io_x[9:0] ? px_buffer_214_g : _GEN_2133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2135 = 10'hd7 == io_x[9:0] ? px_buffer_215_g : _GEN_2134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2136 = 10'hd8 == io_x[9:0] ? px_buffer_216_g : _GEN_2135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2137 = 10'hd9 == io_x[9:0] ? px_buffer_217_g : _GEN_2136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2138 = 10'hda == io_x[9:0] ? px_buffer_218_g : _GEN_2137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2139 = 10'hdb == io_x[9:0] ? px_buffer_219_g : _GEN_2138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2140 = 10'hdc == io_x[9:0] ? px_buffer_220_g : _GEN_2139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2141 = 10'hdd == io_x[9:0] ? px_buffer_221_g : _GEN_2140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2142 = 10'hde == io_x[9:0] ? px_buffer_222_g : _GEN_2141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2143 = 10'hdf == io_x[9:0] ? px_buffer_223_g : _GEN_2142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2144 = 10'he0 == io_x[9:0] ? px_buffer_224_g : _GEN_2143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2145 = 10'he1 == io_x[9:0] ? px_buffer_225_g : _GEN_2144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2146 = 10'he2 == io_x[9:0] ? px_buffer_226_g : _GEN_2145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2147 = 10'he3 == io_x[9:0] ? px_buffer_227_g : _GEN_2146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2148 = 10'he4 == io_x[9:0] ? px_buffer_228_g : _GEN_2147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2149 = 10'he5 == io_x[9:0] ? px_buffer_229_g : _GEN_2148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2150 = 10'he6 == io_x[9:0] ? px_buffer_230_g : _GEN_2149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2151 = 10'he7 == io_x[9:0] ? px_buffer_231_g : _GEN_2150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2152 = 10'he8 == io_x[9:0] ? px_buffer_232_g : _GEN_2151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2153 = 10'he9 == io_x[9:0] ? px_buffer_233_g : _GEN_2152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2154 = 10'hea == io_x[9:0] ? px_buffer_234_g : _GEN_2153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2155 = 10'heb == io_x[9:0] ? px_buffer_235_g : _GEN_2154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2156 = 10'hec == io_x[9:0] ? px_buffer_236_g : _GEN_2155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2157 = 10'hed == io_x[9:0] ? px_buffer_237_g : _GEN_2156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2158 = 10'hee == io_x[9:0] ? px_buffer_238_g : _GEN_2157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2159 = 10'hef == io_x[9:0] ? px_buffer_239_g : _GEN_2158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2160 = 10'hf0 == io_x[9:0] ? px_buffer_240_g : _GEN_2159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2161 = 10'hf1 == io_x[9:0] ? px_buffer_241_g : _GEN_2160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2162 = 10'hf2 == io_x[9:0] ? px_buffer_242_g : _GEN_2161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2163 = 10'hf3 == io_x[9:0] ? px_buffer_243_g : _GEN_2162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2164 = 10'hf4 == io_x[9:0] ? px_buffer_244_g : _GEN_2163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2165 = 10'hf5 == io_x[9:0] ? px_buffer_245_g : _GEN_2164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2166 = 10'hf6 == io_x[9:0] ? px_buffer_246_g : _GEN_2165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2167 = 10'hf7 == io_x[9:0] ? px_buffer_247_g : _GEN_2166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2168 = 10'hf8 == io_x[9:0] ? px_buffer_248_g : _GEN_2167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2169 = 10'hf9 == io_x[9:0] ? px_buffer_249_g : _GEN_2168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2170 = 10'hfa == io_x[9:0] ? px_buffer_250_g : _GEN_2169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2171 = 10'hfb == io_x[9:0] ? px_buffer_251_g : _GEN_2170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2172 = 10'hfc == io_x[9:0] ? px_buffer_252_g : _GEN_2171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2173 = 10'hfd == io_x[9:0] ? px_buffer_253_g : _GEN_2172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2174 = 10'hfe == io_x[9:0] ? px_buffer_254_g : _GEN_2173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2175 = 10'hff == io_x[9:0] ? px_buffer_255_g : _GEN_2174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2176 = 10'h100 == io_x[9:0] ? px_buffer_256_g : _GEN_2175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2177 = 10'h101 == io_x[9:0] ? px_buffer_257_g : _GEN_2176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2178 = 10'h102 == io_x[9:0] ? px_buffer_258_g : _GEN_2177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2179 = 10'h103 == io_x[9:0] ? px_buffer_259_g : _GEN_2178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2180 = 10'h104 == io_x[9:0] ? px_buffer_260_g : _GEN_2179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2181 = 10'h105 == io_x[9:0] ? px_buffer_261_g : _GEN_2180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2182 = 10'h106 == io_x[9:0] ? px_buffer_262_g : _GEN_2181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2183 = 10'h107 == io_x[9:0] ? px_buffer_263_g : _GEN_2182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2184 = 10'h108 == io_x[9:0] ? px_buffer_264_g : _GEN_2183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2185 = 10'h109 == io_x[9:0] ? px_buffer_265_g : _GEN_2184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2186 = 10'h10a == io_x[9:0] ? px_buffer_266_g : _GEN_2185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2187 = 10'h10b == io_x[9:0] ? px_buffer_267_g : _GEN_2186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2188 = 10'h10c == io_x[9:0] ? px_buffer_268_g : _GEN_2187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2189 = 10'h10d == io_x[9:0] ? px_buffer_269_g : _GEN_2188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2190 = 10'h10e == io_x[9:0] ? px_buffer_270_g : _GEN_2189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2191 = 10'h10f == io_x[9:0] ? px_buffer_271_g : _GEN_2190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2192 = 10'h110 == io_x[9:0] ? px_buffer_272_g : _GEN_2191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2193 = 10'h111 == io_x[9:0] ? px_buffer_273_g : _GEN_2192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2194 = 10'h112 == io_x[9:0] ? px_buffer_274_g : _GEN_2193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2195 = 10'h113 == io_x[9:0] ? px_buffer_275_g : _GEN_2194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2196 = 10'h114 == io_x[9:0] ? px_buffer_276_g : _GEN_2195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2197 = 10'h115 == io_x[9:0] ? px_buffer_277_g : _GEN_2196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2198 = 10'h116 == io_x[9:0] ? px_buffer_278_g : _GEN_2197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2199 = 10'h117 == io_x[9:0] ? px_buffer_279_g : _GEN_2198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2200 = 10'h118 == io_x[9:0] ? px_buffer_280_g : _GEN_2199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2201 = 10'h119 == io_x[9:0] ? px_buffer_281_g : _GEN_2200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2202 = 10'h11a == io_x[9:0] ? px_buffer_282_g : _GEN_2201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2203 = 10'h11b == io_x[9:0] ? px_buffer_283_g : _GEN_2202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2204 = 10'h11c == io_x[9:0] ? px_buffer_284_g : _GEN_2203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2205 = 10'h11d == io_x[9:0] ? px_buffer_285_g : _GEN_2204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2206 = 10'h11e == io_x[9:0] ? px_buffer_286_g : _GEN_2205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2207 = 10'h11f == io_x[9:0] ? px_buffer_287_g : _GEN_2206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2208 = 10'h120 == io_x[9:0] ? px_buffer_288_g : _GEN_2207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2209 = 10'h121 == io_x[9:0] ? px_buffer_289_g : _GEN_2208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2210 = 10'h122 == io_x[9:0] ? px_buffer_290_g : _GEN_2209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2211 = 10'h123 == io_x[9:0] ? px_buffer_291_g : _GEN_2210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2212 = 10'h124 == io_x[9:0] ? px_buffer_292_g : _GEN_2211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2213 = 10'h125 == io_x[9:0] ? px_buffer_293_g : _GEN_2212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2214 = 10'h126 == io_x[9:0] ? px_buffer_294_g : _GEN_2213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2215 = 10'h127 == io_x[9:0] ? px_buffer_295_g : _GEN_2214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2216 = 10'h128 == io_x[9:0] ? px_buffer_296_g : _GEN_2215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2217 = 10'h129 == io_x[9:0] ? px_buffer_297_g : _GEN_2216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2218 = 10'h12a == io_x[9:0] ? px_buffer_298_g : _GEN_2217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2219 = 10'h12b == io_x[9:0] ? px_buffer_299_g : _GEN_2218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2220 = 10'h12c == io_x[9:0] ? px_buffer_300_g : _GEN_2219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2221 = 10'h12d == io_x[9:0] ? px_buffer_301_g : _GEN_2220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2222 = 10'h12e == io_x[9:0] ? px_buffer_302_g : _GEN_2221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2223 = 10'h12f == io_x[9:0] ? px_buffer_303_g : _GEN_2222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2224 = 10'h130 == io_x[9:0] ? px_buffer_304_g : _GEN_2223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2225 = 10'h131 == io_x[9:0] ? px_buffer_305_g : _GEN_2224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2226 = 10'h132 == io_x[9:0] ? px_buffer_306_g : _GEN_2225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2227 = 10'h133 == io_x[9:0] ? px_buffer_307_g : _GEN_2226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2228 = 10'h134 == io_x[9:0] ? px_buffer_308_g : _GEN_2227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2229 = 10'h135 == io_x[9:0] ? px_buffer_309_g : _GEN_2228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2230 = 10'h136 == io_x[9:0] ? px_buffer_310_g : _GEN_2229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2231 = 10'h137 == io_x[9:0] ? px_buffer_311_g : _GEN_2230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2232 = 10'h138 == io_x[9:0] ? px_buffer_312_g : _GEN_2231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2233 = 10'h139 == io_x[9:0] ? px_buffer_313_g : _GEN_2232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2234 = 10'h13a == io_x[9:0] ? px_buffer_314_g : _GEN_2233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2235 = 10'h13b == io_x[9:0] ? px_buffer_315_g : _GEN_2234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2236 = 10'h13c == io_x[9:0] ? px_buffer_316_g : _GEN_2235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2237 = 10'h13d == io_x[9:0] ? px_buffer_317_g : _GEN_2236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2238 = 10'h13e == io_x[9:0] ? px_buffer_318_g : _GEN_2237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2239 = 10'h13f == io_x[9:0] ? px_buffer_319_g : _GEN_2238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2240 = 10'h140 == io_x[9:0] ? px_buffer_320_g : _GEN_2239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2241 = 10'h141 == io_x[9:0] ? px_buffer_321_g : _GEN_2240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2242 = 10'h142 == io_x[9:0] ? px_buffer_322_g : _GEN_2241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2243 = 10'h143 == io_x[9:0] ? px_buffer_323_g : _GEN_2242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2244 = 10'h144 == io_x[9:0] ? px_buffer_324_g : _GEN_2243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2245 = 10'h145 == io_x[9:0] ? px_buffer_325_g : _GEN_2244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2246 = 10'h146 == io_x[9:0] ? px_buffer_326_g : _GEN_2245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2247 = 10'h147 == io_x[9:0] ? px_buffer_327_g : _GEN_2246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2248 = 10'h148 == io_x[9:0] ? px_buffer_328_g : _GEN_2247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2249 = 10'h149 == io_x[9:0] ? px_buffer_329_g : _GEN_2248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2250 = 10'h14a == io_x[9:0] ? px_buffer_330_g : _GEN_2249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2251 = 10'h14b == io_x[9:0] ? px_buffer_331_g : _GEN_2250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2252 = 10'h14c == io_x[9:0] ? px_buffer_332_g : _GEN_2251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2253 = 10'h14d == io_x[9:0] ? px_buffer_333_g : _GEN_2252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2254 = 10'h14e == io_x[9:0] ? px_buffer_334_g : _GEN_2253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2255 = 10'h14f == io_x[9:0] ? px_buffer_335_g : _GEN_2254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2256 = 10'h150 == io_x[9:0] ? px_buffer_336_g : _GEN_2255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2257 = 10'h151 == io_x[9:0] ? px_buffer_337_g : _GEN_2256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2258 = 10'h152 == io_x[9:0] ? px_buffer_338_g : _GEN_2257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2259 = 10'h153 == io_x[9:0] ? px_buffer_339_g : _GEN_2258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2260 = 10'h154 == io_x[9:0] ? px_buffer_340_g : _GEN_2259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2261 = 10'h155 == io_x[9:0] ? px_buffer_341_g : _GEN_2260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2262 = 10'h156 == io_x[9:0] ? px_buffer_342_g : _GEN_2261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2263 = 10'h157 == io_x[9:0] ? px_buffer_343_g : _GEN_2262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2264 = 10'h158 == io_x[9:0] ? px_buffer_344_g : _GEN_2263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2265 = 10'h159 == io_x[9:0] ? px_buffer_345_g : _GEN_2264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2266 = 10'h15a == io_x[9:0] ? px_buffer_346_g : _GEN_2265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2267 = 10'h15b == io_x[9:0] ? px_buffer_347_g : _GEN_2266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2268 = 10'h15c == io_x[9:0] ? px_buffer_348_g : _GEN_2267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2269 = 10'h15d == io_x[9:0] ? px_buffer_349_g : _GEN_2268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2270 = 10'h15e == io_x[9:0] ? px_buffer_350_g : _GEN_2269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2271 = 10'h15f == io_x[9:0] ? px_buffer_351_g : _GEN_2270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2272 = 10'h160 == io_x[9:0] ? px_buffer_352_g : _GEN_2271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2273 = 10'h161 == io_x[9:0] ? px_buffer_353_g : _GEN_2272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2274 = 10'h162 == io_x[9:0] ? px_buffer_354_g : _GEN_2273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2275 = 10'h163 == io_x[9:0] ? px_buffer_355_g : _GEN_2274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2276 = 10'h164 == io_x[9:0] ? px_buffer_356_g : _GEN_2275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2277 = 10'h165 == io_x[9:0] ? px_buffer_357_g : _GEN_2276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2278 = 10'h166 == io_x[9:0] ? px_buffer_358_g : _GEN_2277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2279 = 10'h167 == io_x[9:0] ? px_buffer_359_g : _GEN_2278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2280 = 10'h168 == io_x[9:0] ? px_buffer_360_g : _GEN_2279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2281 = 10'h169 == io_x[9:0] ? px_buffer_361_g : _GEN_2280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2282 = 10'h16a == io_x[9:0] ? px_buffer_362_g : _GEN_2281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2283 = 10'h16b == io_x[9:0] ? px_buffer_363_g : _GEN_2282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2284 = 10'h16c == io_x[9:0] ? px_buffer_364_g : _GEN_2283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2285 = 10'h16d == io_x[9:0] ? px_buffer_365_g : _GEN_2284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2286 = 10'h16e == io_x[9:0] ? px_buffer_366_g : _GEN_2285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2287 = 10'h16f == io_x[9:0] ? px_buffer_367_g : _GEN_2286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2288 = 10'h170 == io_x[9:0] ? px_buffer_368_g : _GEN_2287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2289 = 10'h171 == io_x[9:0] ? px_buffer_369_g : _GEN_2288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2290 = 10'h172 == io_x[9:0] ? px_buffer_370_g : _GEN_2289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2291 = 10'h173 == io_x[9:0] ? px_buffer_371_g : _GEN_2290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2292 = 10'h174 == io_x[9:0] ? px_buffer_372_g : _GEN_2291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2293 = 10'h175 == io_x[9:0] ? px_buffer_373_g : _GEN_2292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2294 = 10'h176 == io_x[9:0] ? px_buffer_374_g : _GEN_2293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2295 = 10'h177 == io_x[9:0] ? px_buffer_375_g : _GEN_2294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2296 = 10'h178 == io_x[9:0] ? px_buffer_376_g : _GEN_2295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2297 = 10'h179 == io_x[9:0] ? px_buffer_377_g : _GEN_2296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2298 = 10'h17a == io_x[9:0] ? px_buffer_378_g : _GEN_2297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2299 = 10'h17b == io_x[9:0] ? px_buffer_379_g : _GEN_2298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2300 = 10'h17c == io_x[9:0] ? px_buffer_380_g : _GEN_2299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2301 = 10'h17d == io_x[9:0] ? px_buffer_381_g : _GEN_2300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2302 = 10'h17e == io_x[9:0] ? px_buffer_382_g : _GEN_2301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2303 = 10'h17f == io_x[9:0] ? px_buffer_383_g : _GEN_2302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2304 = 10'h180 == io_x[9:0] ? px_buffer_384_g : _GEN_2303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2305 = 10'h181 == io_x[9:0] ? px_buffer_385_g : _GEN_2304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2306 = 10'h182 == io_x[9:0] ? px_buffer_386_g : _GEN_2305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2307 = 10'h183 == io_x[9:0] ? px_buffer_387_g : _GEN_2306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2308 = 10'h184 == io_x[9:0] ? px_buffer_388_g : _GEN_2307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2309 = 10'h185 == io_x[9:0] ? px_buffer_389_g : _GEN_2308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2310 = 10'h186 == io_x[9:0] ? px_buffer_390_g : _GEN_2309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2311 = 10'h187 == io_x[9:0] ? px_buffer_391_g : _GEN_2310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2312 = 10'h188 == io_x[9:0] ? px_buffer_392_g : _GEN_2311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2313 = 10'h189 == io_x[9:0] ? px_buffer_393_g : _GEN_2312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2314 = 10'h18a == io_x[9:0] ? px_buffer_394_g : _GEN_2313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2315 = 10'h18b == io_x[9:0] ? px_buffer_395_g : _GEN_2314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2316 = 10'h18c == io_x[9:0] ? px_buffer_396_g : _GEN_2315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2317 = 10'h18d == io_x[9:0] ? px_buffer_397_g : _GEN_2316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2318 = 10'h18e == io_x[9:0] ? px_buffer_398_g : _GEN_2317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2319 = 10'h18f == io_x[9:0] ? px_buffer_399_g : _GEN_2318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2320 = 10'h190 == io_x[9:0] ? px_buffer_400_g : _GEN_2319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2321 = 10'h191 == io_x[9:0] ? px_buffer_401_g : _GEN_2320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2322 = 10'h192 == io_x[9:0] ? px_buffer_402_g : _GEN_2321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2323 = 10'h193 == io_x[9:0] ? px_buffer_403_g : _GEN_2322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2324 = 10'h194 == io_x[9:0] ? px_buffer_404_g : _GEN_2323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2325 = 10'h195 == io_x[9:0] ? px_buffer_405_g : _GEN_2324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2326 = 10'h196 == io_x[9:0] ? px_buffer_406_g : _GEN_2325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2327 = 10'h197 == io_x[9:0] ? px_buffer_407_g : _GEN_2326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2328 = 10'h198 == io_x[9:0] ? px_buffer_408_g : _GEN_2327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2329 = 10'h199 == io_x[9:0] ? px_buffer_409_g : _GEN_2328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2330 = 10'h19a == io_x[9:0] ? px_buffer_410_g : _GEN_2329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2331 = 10'h19b == io_x[9:0] ? px_buffer_411_g : _GEN_2330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2332 = 10'h19c == io_x[9:0] ? px_buffer_412_g : _GEN_2331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2333 = 10'h19d == io_x[9:0] ? px_buffer_413_g : _GEN_2332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2334 = 10'h19e == io_x[9:0] ? px_buffer_414_g : _GEN_2333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2335 = 10'h19f == io_x[9:0] ? px_buffer_415_g : _GEN_2334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2336 = 10'h1a0 == io_x[9:0] ? px_buffer_416_g : _GEN_2335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2337 = 10'h1a1 == io_x[9:0] ? px_buffer_417_g : _GEN_2336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2338 = 10'h1a2 == io_x[9:0] ? px_buffer_418_g : _GEN_2337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2339 = 10'h1a3 == io_x[9:0] ? px_buffer_419_g : _GEN_2338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2340 = 10'h1a4 == io_x[9:0] ? px_buffer_420_g : _GEN_2339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2341 = 10'h1a5 == io_x[9:0] ? px_buffer_421_g : _GEN_2340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2342 = 10'h1a6 == io_x[9:0] ? px_buffer_422_g : _GEN_2341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2343 = 10'h1a7 == io_x[9:0] ? px_buffer_423_g : _GEN_2342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2344 = 10'h1a8 == io_x[9:0] ? px_buffer_424_g : _GEN_2343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2345 = 10'h1a9 == io_x[9:0] ? px_buffer_425_g : _GEN_2344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2346 = 10'h1aa == io_x[9:0] ? px_buffer_426_g : _GEN_2345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2347 = 10'h1ab == io_x[9:0] ? px_buffer_427_g : _GEN_2346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2348 = 10'h1ac == io_x[9:0] ? px_buffer_428_g : _GEN_2347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2349 = 10'h1ad == io_x[9:0] ? px_buffer_429_g : _GEN_2348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2350 = 10'h1ae == io_x[9:0] ? px_buffer_430_g : _GEN_2349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2351 = 10'h1af == io_x[9:0] ? px_buffer_431_g : _GEN_2350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2352 = 10'h1b0 == io_x[9:0] ? px_buffer_432_g : _GEN_2351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2353 = 10'h1b1 == io_x[9:0] ? px_buffer_433_g : _GEN_2352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2354 = 10'h1b2 == io_x[9:0] ? px_buffer_434_g : _GEN_2353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2355 = 10'h1b3 == io_x[9:0] ? px_buffer_435_g : _GEN_2354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2356 = 10'h1b4 == io_x[9:0] ? px_buffer_436_g : _GEN_2355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2357 = 10'h1b5 == io_x[9:0] ? px_buffer_437_g : _GEN_2356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2358 = 10'h1b6 == io_x[9:0] ? px_buffer_438_g : _GEN_2357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2359 = 10'h1b7 == io_x[9:0] ? px_buffer_439_g : _GEN_2358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2360 = 10'h1b8 == io_x[9:0] ? px_buffer_440_g : _GEN_2359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2361 = 10'h1b9 == io_x[9:0] ? px_buffer_441_g : _GEN_2360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2362 = 10'h1ba == io_x[9:0] ? px_buffer_442_g : _GEN_2361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2363 = 10'h1bb == io_x[9:0] ? px_buffer_443_g : _GEN_2362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2364 = 10'h1bc == io_x[9:0] ? px_buffer_444_g : _GEN_2363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2365 = 10'h1bd == io_x[9:0] ? px_buffer_445_g : _GEN_2364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2366 = 10'h1be == io_x[9:0] ? px_buffer_446_g : _GEN_2365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2367 = 10'h1bf == io_x[9:0] ? px_buffer_447_g : _GEN_2366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2368 = 10'h1c0 == io_x[9:0] ? px_buffer_448_g : _GEN_2367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2369 = 10'h1c1 == io_x[9:0] ? px_buffer_449_g : _GEN_2368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2370 = 10'h1c2 == io_x[9:0] ? px_buffer_450_g : _GEN_2369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2371 = 10'h1c3 == io_x[9:0] ? px_buffer_451_g : _GEN_2370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2372 = 10'h1c4 == io_x[9:0] ? px_buffer_452_g : _GEN_2371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2373 = 10'h1c5 == io_x[9:0] ? px_buffer_453_g : _GEN_2372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2374 = 10'h1c6 == io_x[9:0] ? px_buffer_454_g : _GEN_2373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2375 = 10'h1c7 == io_x[9:0] ? px_buffer_455_g : _GEN_2374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2376 = 10'h1c8 == io_x[9:0] ? px_buffer_456_g : _GEN_2375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2377 = 10'h1c9 == io_x[9:0] ? px_buffer_457_g : _GEN_2376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2378 = 10'h1ca == io_x[9:0] ? px_buffer_458_g : _GEN_2377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2379 = 10'h1cb == io_x[9:0] ? px_buffer_459_g : _GEN_2378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2380 = 10'h1cc == io_x[9:0] ? px_buffer_460_g : _GEN_2379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2381 = 10'h1cd == io_x[9:0] ? px_buffer_461_g : _GEN_2380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2382 = 10'h1ce == io_x[9:0] ? px_buffer_462_g : _GEN_2381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2383 = 10'h1cf == io_x[9:0] ? px_buffer_463_g : _GEN_2382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2384 = 10'h1d0 == io_x[9:0] ? px_buffer_464_g : _GEN_2383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2385 = 10'h1d1 == io_x[9:0] ? px_buffer_465_g : _GEN_2384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2386 = 10'h1d2 == io_x[9:0] ? px_buffer_466_g : _GEN_2385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2387 = 10'h1d3 == io_x[9:0] ? px_buffer_467_g : _GEN_2386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2388 = 10'h1d4 == io_x[9:0] ? px_buffer_468_g : _GEN_2387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2389 = 10'h1d5 == io_x[9:0] ? px_buffer_469_g : _GEN_2388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2390 = 10'h1d6 == io_x[9:0] ? px_buffer_470_g : _GEN_2389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2391 = 10'h1d7 == io_x[9:0] ? px_buffer_471_g : _GEN_2390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2392 = 10'h1d8 == io_x[9:0] ? px_buffer_472_g : _GEN_2391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2393 = 10'h1d9 == io_x[9:0] ? px_buffer_473_g : _GEN_2392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2394 = 10'h1da == io_x[9:0] ? px_buffer_474_g : _GEN_2393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2395 = 10'h1db == io_x[9:0] ? px_buffer_475_g : _GEN_2394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2396 = 10'h1dc == io_x[9:0] ? px_buffer_476_g : _GEN_2395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2397 = 10'h1dd == io_x[9:0] ? px_buffer_477_g : _GEN_2396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2398 = 10'h1de == io_x[9:0] ? px_buffer_478_g : _GEN_2397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2399 = 10'h1df == io_x[9:0] ? px_buffer_479_g : _GEN_2398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2400 = 10'h1e0 == io_x[9:0] ? px_buffer_480_g : _GEN_2399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2401 = 10'h1e1 == io_x[9:0] ? px_buffer_481_g : _GEN_2400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2402 = 10'h1e2 == io_x[9:0] ? px_buffer_482_g : _GEN_2401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2403 = 10'h1e3 == io_x[9:0] ? px_buffer_483_g : _GEN_2402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2404 = 10'h1e4 == io_x[9:0] ? px_buffer_484_g : _GEN_2403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2405 = 10'h1e5 == io_x[9:0] ? px_buffer_485_g : _GEN_2404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2406 = 10'h1e6 == io_x[9:0] ? px_buffer_486_g : _GEN_2405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2407 = 10'h1e7 == io_x[9:0] ? px_buffer_487_g : _GEN_2406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2408 = 10'h1e8 == io_x[9:0] ? px_buffer_488_g : _GEN_2407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2409 = 10'h1e9 == io_x[9:0] ? px_buffer_489_g : _GEN_2408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2410 = 10'h1ea == io_x[9:0] ? px_buffer_490_g : _GEN_2409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2411 = 10'h1eb == io_x[9:0] ? px_buffer_491_g : _GEN_2410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2412 = 10'h1ec == io_x[9:0] ? px_buffer_492_g : _GEN_2411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2413 = 10'h1ed == io_x[9:0] ? px_buffer_493_g : _GEN_2412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2414 = 10'h1ee == io_x[9:0] ? px_buffer_494_g : _GEN_2413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2415 = 10'h1ef == io_x[9:0] ? px_buffer_495_g : _GEN_2414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2416 = 10'h1f0 == io_x[9:0] ? px_buffer_496_g : _GEN_2415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2417 = 10'h1f1 == io_x[9:0] ? px_buffer_497_g : _GEN_2416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2418 = 10'h1f2 == io_x[9:0] ? px_buffer_498_g : _GEN_2417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2419 = 10'h1f3 == io_x[9:0] ? px_buffer_499_g : _GEN_2418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2420 = 10'h1f4 == io_x[9:0] ? px_buffer_500_g : _GEN_2419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2421 = 10'h1f5 == io_x[9:0] ? px_buffer_501_g : _GEN_2420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2422 = 10'h1f6 == io_x[9:0] ? px_buffer_502_g : _GEN_2421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2423 = 10'h1f7 == io_x[9:0] ? px_buffer_503_g : _GEN_2422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2424 = 10'h1f8 == io_x[9:0] ? px_buffer_504_g : _GEN_2423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2425 = 10'h1f9 == io_x[9:0] ? px_buffer_505_g : _GEN_2424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2426 = 10'h1fa == io_x[9:0] ? px_buffer_506_g : _GEN_2425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2427 = 10'h1fb == io_x[9:0] ? px_buffer_507_g : _GEN_2426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2428 = 10'h1fc == io_x[9:0] ? px_buffer_508_g : _GEN_2427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2429 = 10'h1fd == io_x[9:0] ? px_buffer_509_g : _GEN_2428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2430 = 10'h1fe == io_x[9:0] ? px_buffer_510_g : _GEN_2429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2431 = 10'h1ff == io_x[9:0] ? px_buffer_511_g : _GEN_2430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2432 = 10'h200 == io_x[9:0] ? px_buffer_512_g : _GEN_2431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2433 = 10'h201 == io_x[9:0] ? px_buffer_513_g : _GEN_2432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2434 = 10'h202 == io_x[9:0] ? px_buffer_514_g : _GEN_2433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2435 = 10'h203 == io_x[9:0] ? px_buffer_515_g : _GEN_2434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2436 = 10'h204 == io_x[9:0] ? px_buffer_516_g : _GEN_2435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2437 = 10'h205 == io_x[9:0] ? px_buffer_517_g : _GEN_2436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2438 = 10'h206 == io_x[9:0] ? px_buffer_518_g : _GEN_2437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2439 = 10'h207 == io_x[9:0] ? px_buffer_519_g : _GEN_2438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2440 = 10'h208 == io_x[9:0] ? px_buffer_520_g : _GEN_2439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2441 = 10'h209 == io_x[9:0] ? px_buffer_521_g : _GEN_2440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2442 = 10'h20a == io_x[9:0] ? px_buffer_522_g : _GEN_2441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2443 = 10'h20b == io_x[9:0] ? px_buffer_523_g : _GEN_2442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2444 = 10'h20c == io_x[9:0] ? px_buffer_524_g : _GEN_2443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2445 = 10'h20d == io_x[9:0] ? px_buffer_525_g : _GEN_2444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2446 = 10'h20e == io_x[9:0] ? px_buffer_526_g : _GEN_2445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2447 = 10'h20f == io_x[9:0] ? px_buffer_527_g : _GEN_2446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2448 = 10'h210 == io_x[9:0] ? px_buffer_528_g : _GEN_2447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2449 = 10'h211 == io_x[9:0] ? px_buffer_529_g : _GEN_2448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2450 = 10'h212 == io_x[9:0] ? px_buffer_530_g : _GEN_2449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2451 = 10'h213 == io_x[9:0] ? px_buffer_531_g : _GEN_2450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2452 = 10'h214 == io_x[9:0] ? px_buffer_532_g : _GEN_2451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2453 = 10'h215 == io_x[9:0] ? px_buffer_533_g : _GEN_2452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2454 = 10'h216 == io_x[9:0] ? px_buffer_534_g : _GEN_2453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2455 = 10'h217 == io_x[9:0] ? px_buffer_535_g : _GEN_2454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2456 = 10'h218 == io_x[9:0] ? px_buffer_536_g : _GEN_2455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2457 = 10'h219 == io_x[9:0] ? px_buffer_537_g : _GEN_2456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2458 = 10'h21a == io_x[9:0] ? px_buffer_538_g : _GEN_2457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2459 = 10'h21b == io_x[9:0] ? px_buffer_539_g : _GEN_2458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2460 = 10'h21c == io_x[9:0] ? px_buffer_540_g : _GEN_2459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2461 = 10'h21d == io_x[9:0] ? px_buffer_541_g : _GEN_2460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2462 = 10'h21e == io_x[9:0] ? px_buffer_542_g : _GEN_2461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2463 = 10'h21f == io_x[9:0] ? px_buffer_543_g : _GEN_2462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2464 = 10'h220 == io_x[9:0] ? px_buffer_544_g : _GEN_2463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2465 = 10'h221 == io_x[9:0] ? px_buffer_545_g : _GEN_2464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2466 = 10'h222 == io_x[9:0] ? px_buffer_546_g : _GEN_2465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2467 = 10'h223 == io_x[9:0] ? px_buffer_547_g : _GEN_2466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2468 = 10'h224 == io_x[9:0] ? px_buffer_548_g : _GEN_2467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2469 = 10'h225 == io_x[9:0] ? px_buffer_549_g : _GEN_2468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2470 = 10'h226 == io_x[9:0] ? px_buffer_550_g : _GEN_2469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2471 = 10'h227 == io_x[9:0] ? px_buffer_551_g : _GEN_2470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2472 = 10'h228 == io_x[9:0] ? px_buffer_552_g : _GEN_2471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2473 = 10'h229 == io_x[9:0] ? px_buffer_553_g : _GEN_2472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2474 = 10'h22a == io_x[9:0] ? px_buffer_554_g : _GEN_2473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2475 = 10'h22b == io_x[9:0] ? px_buffer_555_g : _GEN_2474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2476 = 10'h22c == io_x[9:0] ? px_buffer_556_g : _GEN_2475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2477 = 10'h22d == io_x[9:0] ? px_buffer_557_g : _GEN_2476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2478 = 10'h22e == io_x[9:0] ? px_buffer_558_g : _GEN_2477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2479 = 10'h22f == io_x[9:0] ? px_buffer_559_g : _GEN_2478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2480 = 10'h230 == io_x[9:0] ? px_buffer_560_g : _GEN_2479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2481 = 10'h231 == io_x[9:0] ? px_buffer_561_g : _GEN_2480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2482 = 10'h232 == io_x[9:0] ? px_buffer_562_g : _GEN_2481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2483 = 10'h233 == io_x[9:0] ? px_buffer_563_g : _GEN_2482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2484 = 10'h234 == io_x[9:0] ? px_buffer_564_g : _GEN_2483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2485 = 10'h235 == io_x[9:0] ? px_buffer_565_g : _GEN_2484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2486 = 10'h236 == io_x[9:0] ? px_buffer_566_g : _GEN_2485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2487 = 10'h237 == io_x[9:0] ? px_buffer_567_g : _GEN_2486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2488 = 10'h238 == io_x[9:0] ? px_buffer_568_g : _GEN_2487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2489 = 10'h239 == io_x[9:0] ? px_buffer_569_g : _GEN_2488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2490 = 10'h23a == io_x[9:0] ? px_buffer_570_g : _GEN_2489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2491 = 10'h23b == io_x[9:0] ? px_buffer_571_g : _GEN_2490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2492 = 10'h23c == io_x[9:0] ? px_buffer_572_g : _GEN_2491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2493 = 10'h23d == io_x[9:0] ? px_buffer_573_g : _GEN_2492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2494 = 10'h23e == io_x[9:0] ? px_buffer_574_g : _GEN_2493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2495 = 10'h23f == io_x[9:0] ? px_buffer_575_g : _GEN_2494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2496 = 10'h240 == io_x[9:0] ? px_buffer_576_g : _GEN_2495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2497 = 10'h241 == io_x[9:0] ? px_buffer_577_g : _GEN_2496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2498 = 10'h242 == io_x[9:0] ? px_buffer_578_g : _GEN_2497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2499 = 10'h243 == io_x[9:0] ? px_buffer_579_g : _GEN_2498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2500 = 10'h244 == io_x[9:0] ? px_buffer_580_g : _GEN_2499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2501 = 10'h245 == io_x[9:0] ? px_buffer_581_g : _GEN_2500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2502 = 10'h246 == io_x[9:0] ? px_buffer_582_g : _GEN_2501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2503 = 10'h247 == io_x[9:0] ? px_buffer_583_g : _GEN_2502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2504 = 10'h248 == io_x[9:0] ? px_buffer_584_g : _GEN_2503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2505 = 10'h249 == io_x[9:0] ? px_buffer_585_g : _GEN_2504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2506 = 10'h24a == io_x[9:0] ? px_buffer_586_g : _GEN_2505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2507 = 10'h24b == io_x[9:0] ? px_buffer_587_g : _GEN_2506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2508 = 10'h24c == io_x[9:0] ? px_buffer_588_g : _GEN_2507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2509 = 10'h24d == io_x[9:0] ? px_buffer_589_g : _GEN_2508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2510 = 10'h24e == io_x[9:0] ? px_buffer_590_g : _GEN_2509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2511 = 10'h24f == io_x[9:0] ? px_buffer_591_g : _GEN_2510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2512 = 10'h250 == io_x[9:0] ? px_buffer_592_g : _GEN_2511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2513 = 10'h251 == io_x[9:0] ? px_buffer_593_g : _GEN_2512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2514 = 10'h252 == io_x[9:0] ? px_buffer_594_g : _GEN_2513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2515 = 10'h253 == io_x[9:0] ? px_buffer_595_g : _GEN_2514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2516 = 10'h254 == io_x[9:0] ? px_buffer_596_g : _GEN_2515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2517 = 10'h255 == io_x[9:0] ? px_buffer_597_g : _GEN_2516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2518 = 10'h256 == io_x[9:0] ? px_buffer_598_g : _GEN_2517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2519 = 10'h257 == io_x[9:0] ? px_buffer_599_g : _GEN_2518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2520 = 10'h258 == io_x[9:0] ? px_buffer_600_g : _GEN_2519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2521 = 10'h259 == io_x[9:0] ? px_buffer_601_g : _GEN_2520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2522 = 10'h25a == io_x[9:0] ? px_buffer_602_g : _GEN_2521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2523 = 10'h25b == io_x[9:0] ? px_buffer_603_g : _GEN_2522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2524 = 10'h25c == io_x[9:0] ? px_buffer_604_g : _GEN_2523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2525 = 10'h25d == io_x[9:0] ? px_buffer_605_g : _GEN_2524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2526 = 10'h25e == io_x[9:0] ? px_buffer_606_g : _GEN_2525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2527 = 10'h25f == io_x[9:0] ? px_buffer_607_g : _GEN_2526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2528 = 10'h260 == io_x[9:0] ? px_buffer_608_g : _GEN_2527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2529 = 10'h261 == io_x[9:0] ? px_buffer_609_g : _GEN_2528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2530 = 10'h262 == io_x[9:0] ? px_buffer_610_g : _GEN_2529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2531 = 10'h263 == io_x[9:0] ? px_buffer_611_g : _GEN_2530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2532 = 10'h264 == io_x[9:0] ? px_buffer_612_g : _GEN_2531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2533 = 10'h265 == io_x[9:0] ? px_buffer_613_g : _GEN_2532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2534 = 10'h266 == io_x[9:0] ? px_buffer_614_g : _GEN_2533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2535 = 10'h267 == io_x[9:0] ? px_buffer_615_g : _GEN_2534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2536 = 10'h268 == io_x[9:0] ? px_buffer_616_g : _GEN_2535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2537 = 10'h269 == io_x[9:0] ? px_buffer_617_g : _GEN_2536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2538 = 10'h26a == io_x[9:0] ? px_buffer_618_g : _GEN_2537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2539 = 10'h26b == io_x[9:0] ? px_buffer_619_g : _GEN_2538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2540 = 10'h26c == io_x[9:0] ? px_buffer_620_g : _GEN_2539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2541 = 10'h26d == io_x[9:0] ? px_buffer_621_g : _GEN_2540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2542 = 10'h26e == io_x[9:0] ? px_buffer_622_g : _GEN_2541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2543 = 10'h26f == io_x[9:0] ? px_buffer_623_g : _GEN_2542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2544 = 10'h270 == io_x[9:0] ? px_buffer_624_g : _GEN_2543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2545 = 10'h271 == io_x[9:0] ? px_buffer_625_g : _GEN_2544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2546 = 10'h272 == io_x[9:0] ? px_buffer_626_g : _GEN_2545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2547 = 10'h273 == io_x[9:0] ? px_buffer_627_g : _GEN_2546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2548 = 10'h274 == io_x[9:0] ? px_buffer_628_g : _GEN_2547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2549 = 10'h275 == io_x[9:0] ? px_buffer_629_g : _GEN_2548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2550 = 10'h276 == io_x[9:0] ? px_buffer_630_g : _GEN_2549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2551 = 10'h277 == io_x[9:0] ? px_buffer_631_g : _GEN_2550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2552 = 10'h278 == io_x[9:0] ? px_buffer_632_g : _GEN_2551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2553 = 10'h279 == io_x[9:0] ? px_buffer_633_g : _GEN_2552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2554 = 10'h27a == io_x[9:0] ? px_buffer_634_g : _GEN_2553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2555 = 10'h27b == io_x[9:0] ? px_buffer_635_g : _GEN_2554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2556 = 10'h27c == io_x[9:0] ? px_buffer_636_g : _GEN_2555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2557 = 10'h27d == io_x[9:0] ? px_buffer_637_g : _GEN_2556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2558 = 10'h27e == io_x[9:0] ? px_buffer_638_g : _GEN_2557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2559 = 10'h27f == io_x[9:0] ? px_buffer_639_g : _GEN_2558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _T_83 = {1'h0,_GEN_2559}; // @[EdgeDetect.scala 57:47]
  wire [8:0] _T_85 = {1'h0,last_px_g}; // @[EdgeDetect.scala 57:79]
  wire [8:0] _T_88 = $signed(_T_83) - $signed(_T_85); // @[EdgeDetect.scala 57:54]
  assign io_px_out_r = _T_14[8:1]; // @[EdgeDetect.scala 39:36]
  assign io_px_out_g = _T_32[8:1]; // @[EdgeDetect.scala 44:36]
  assign io_px_out_b = _T_32[8:1]; // @[EdgeDetect.scala 44:36]
  always @(posedge clock) begin
    if (10'h0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_0_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_0_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_0_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_0_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_1_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_1_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_1_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_1_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_2_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_2_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_2_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_2_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_3_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_3_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_3_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_3_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_4_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_4_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_4_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_4_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_5_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_5_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_5_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_5_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_6_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_6_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_6_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_6_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_7_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_7_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_7_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_7_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_8_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_8_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_8_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_8_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_9_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_9_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_9_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_9_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_10_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_10_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_10_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_10_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_11_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_11_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_11_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_11_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_12_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_12_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_12_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_12_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_13_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_13_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_13_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_13_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_14_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_14_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_14_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_14_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_15_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_15_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_15_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_15_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_16_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_16_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_16_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_16_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_17_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_17_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_17_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_17_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_18_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_18_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_18_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_18_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_19_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_19_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_19_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_19_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_20_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_20_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_20_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_20_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_21_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_21_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_21_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_21_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_22_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_22_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_22_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_22_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_23_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_23_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_23_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_23_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_24_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_24_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_24_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_24_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_25_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_25_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_25_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_25_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_26_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_26_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_26_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_26_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_27_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_27_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_27_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_27_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_28_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_28_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_28_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_28_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_29_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_29_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_29_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_29_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_30_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_30_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_30_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_30_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_31_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_31_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_31_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_31_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_32_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_32_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_32_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_32_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_33_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_33_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_33_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_33_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_34_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_34_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_34_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_34_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_35_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_35_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_35_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_35_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_36_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_36_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_36_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_36_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_37_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_37_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_37_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_37_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_38_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_38_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_38_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_38_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_39_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_39_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_39_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_39_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h28 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_40_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_40_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h28 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_40_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_40_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h29 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_41_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_41_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h29 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_41_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_41_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_42_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_42_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_42_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_42_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_43_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_43_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_43_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_43_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_44_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_44_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_44_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_44_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_45_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_45_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_45_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_45_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_46_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_46_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_46_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_46_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_47_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_47_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h2f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_47_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_47_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h30 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_48_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_48_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h30 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_48_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_48_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h31 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_49_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_49_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h31 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_49_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_49_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h32 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_50_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_50_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h32 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_50_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_50_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h33 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_51_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_51_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h33 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_51_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_51_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h34 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_52_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_52_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h34 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_52_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_52_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h35 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_53_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_53_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h35 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_53_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_53_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h36 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_54_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_54_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h36 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_54_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_54_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h37 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_55_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_55_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h37 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_55_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_55_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h38 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_56_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_56_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h38 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_56_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_56_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h39 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_57_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_57_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h39 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_57_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_57_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_58_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_58_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_58_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_58_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_59_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_59_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_59_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_59_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_60_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_60_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_60_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_60_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_61_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_61_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_61_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_61_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_62_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_62_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_62_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_62_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_63_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_63_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h3f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_63_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_63_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h40 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_64_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_64_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h40 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_64_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_64_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h41 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_65_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_65_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h41 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_65_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_65_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h42 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_66_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_66_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h42 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_66_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_66_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h43 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_67_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_67_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h43 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_67_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_67_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h44 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_68_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_68_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h44 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_68_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_68_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h45 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_69_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_69_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h45 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_69_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_69_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h46 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_70_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_70_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h46 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_70_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_70_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h47 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_71_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_71_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h47 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_71_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_71_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h48 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_72_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_72_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h48 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_72_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_72_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h49 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_73_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_73_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h49 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_73_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_73_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_74_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_74_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_74_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_74_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_75_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_75_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_75_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_75_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_76_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_76_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_76_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_76_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_77_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_77_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_77_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_77_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_78_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_78_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_78_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_78_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_79_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_79_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h4f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_79_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_79_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h50 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_80_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_80_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h50 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_80_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_80_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h51 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_81_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_81_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h51 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_81_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_81_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h52 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_82_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_82_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h52 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_82_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_82_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h53 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_83_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_83_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h53 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_83_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_83_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h54 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_84_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_84_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h54 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_84_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_84_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h55 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_85_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_85_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h55 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_85_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_85_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h56 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_86_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_86_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h56 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_86_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_86_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h57 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_87_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_87_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h57 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_87_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_87_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h58 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_88_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_88_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h58 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_88_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_88_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h59 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_89_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_89_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h59 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_89_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_89_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_90_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_90_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_90_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_90_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_91_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_91_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_91_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_91_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_92_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_92_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_92_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_92_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_93_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_93_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_93_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_93_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_94_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_94_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_94_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_94_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_95_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_95_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h5f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_95_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_95_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h60 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_96_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_96_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h60 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_96_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_96_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h61 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_97_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_97_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h61 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_97_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_97_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h62 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_98_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_98_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h62 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_98_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_98_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h63 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_99_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_99_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h63 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_99_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_99_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h64 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_100_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_100_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h64 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_100_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_100_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h65 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_101_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_101_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h65 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_101_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_101_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h66 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_102_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_102_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h66 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_102_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_102_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h67 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_103_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_103_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h67 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_103_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_103_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h68 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_104_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_104_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h68 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_104_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_104_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h69 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_105_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_105_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h69 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_105_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_105_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_106_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_106_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_106_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_106_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_107_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_107_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_107_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_107_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_108_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_108_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_108_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_108_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_109_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_109_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_109_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_109_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_110_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_110_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_110_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_110_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_111_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_111_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h6f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_111_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_111_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h70 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_112_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_112_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h70 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_112_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_112_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h71 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_113_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_113_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h71 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_113_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_113_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h72 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_114_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_114_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h72 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_114_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_114_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h73 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_115_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_115_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h73 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_115_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_115_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h74 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_116_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_116_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h74 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_116_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_116_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h75 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_117_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_117_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h75 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_117_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_117_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h76 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_118_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_118_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h76 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_118_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_118_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h77 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_119_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_119_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h77 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_119_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_119_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h78 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_120_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_120_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h78 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_120_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_120_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h79 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_121_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_121_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h79 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_121_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_121_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_122_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_122_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_122_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_122_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_123_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_123_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_123_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_123_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_124_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_124_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_124_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_124_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_125_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_125_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_125_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_125_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_126_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_126_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_126_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_126_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_127_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_127_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h7f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_127_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_127_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h80 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_128_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_128_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h80 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_128_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_128_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h81 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_129_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_129_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h81 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_129_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_129_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h82 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_130_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_130_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h82 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_130_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_130_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h83 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_131_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_131_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h83 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_131_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_131_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h84 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_132_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_132_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h84 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_132_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_132_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h85 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_133_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_133_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h85 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_133_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_133_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h86 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_134_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_134_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h86 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_134_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_134_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h87 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_135_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_135_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h87 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_135_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_135_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h88 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_136_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_136_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h88 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_136_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_136_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h89 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_137_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_137_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h89 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_137_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_137_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_138_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_138_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_138_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_138_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_139_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_139_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_139_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_139_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_140_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_140_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_140_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_140_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_141_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_141_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_141_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_141_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_142_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_142_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_142_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_142_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_143_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_143_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h8f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_143_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_143_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h90 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_144_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_144_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h90 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_144_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_144_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h91 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_145_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_145_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h91 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_145_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_145_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h92 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_146_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_146_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h92 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_146_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_146_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h93 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_147_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_147_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h93 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_147_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_147_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h94 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_148_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_148_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h94 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_148_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_148_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h95 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_149_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_149_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h95 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_149_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_149_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h96 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_150_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_150_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h96 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_150_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_150_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h97 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_151_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_151_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h97 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_151_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_151_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h98 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_152_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_152_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h98 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_152_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_152_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h99 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_153_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_153_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h99 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_153_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_153_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_154_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_154_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_154_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_154_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_155_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_155_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_155_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_155_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_156_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_156_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_156_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_156_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_157_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_157_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_157_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_157_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_158_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_158_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_158_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_158_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_159_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_159_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h9f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_159_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_159_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_160_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_160_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_160_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_160_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_161_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_161_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_161_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_161_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_162_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_162_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_162_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_162_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_163_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_163_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_163_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_163_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_164_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_164_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_164_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_164_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_165_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_165_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_165_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_165_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_166_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_166_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_166_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_166_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_167_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_167_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_167_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_167_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_168_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_168_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_168_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_168_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_169_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_169_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'ha9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_169_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_169_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'haa == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_170_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_170_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'haa == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_170_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_170_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hab == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_171_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_171_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hab == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_171_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_171_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hac == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_172_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_172_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hac == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_172_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_172_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'had == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_173_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_173_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'had == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_173_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_173_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hae == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_174_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_174_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hae == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_174_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_174_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'haf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_175_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_175_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'haf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_175_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_175_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_176_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_176_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_176_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_176_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_177_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_177_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_177_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_177_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_178_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_178_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_178_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_178_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_179_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_179_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_179_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_179_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_180_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_180_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_180_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_180_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_181_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_181_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_181_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_181_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_182_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_182_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_182_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_182_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_183_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_183_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_183_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_183_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_184_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_184_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_184_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_184_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_185_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_185_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hb9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_185_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_185_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hba == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_186_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_186_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hba == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_186_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_186_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_187_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_187_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_187_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_187_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_188_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_188_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_188_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_188_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_189_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_189_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_189_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_189_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbe == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_190_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_190_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbe == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_190_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_190_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_191_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_191_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hbf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_191_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_191_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_192_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_192_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_192_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_192_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_193_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_193_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_193_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_193_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_194_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_194_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_194_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_194_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_195_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_195_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_195_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_195_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_196_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_196_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_196_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_196_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_197_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_197_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_197_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_197_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_198_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_198_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_198_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_198_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_199_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_199_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_199_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_199_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_200_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_200_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_200_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_200_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_201_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_201_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hc9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_201_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_201_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hca == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_202_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_202_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hca == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_202_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_202_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hcb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_203_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_203_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hcb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_203_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_203_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hcc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_204_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_204_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hcc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_204_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_204_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hcd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_205_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_205_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hcd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_205_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_205_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hce == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_206_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_206_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hce == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_206_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_206_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hcf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_207_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_207_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hcf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_207_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_207_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_208_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_208_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_208_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_208_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_209_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_209_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_209_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_209_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_210_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_210_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_210_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_210_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_211_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_211_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_211_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_211_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_212_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_212_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_212_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_212_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_213_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_213_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_213_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_213_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_214_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_214_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_214_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_214_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_215_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_215_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_215_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_215_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_216_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_216_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_216_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_216_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_217_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_217_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hd9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_217_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_217_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hda == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_218_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_218_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hda == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_218_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_218_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hdb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_219_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_219_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hdb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_219_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_219_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hdc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_220_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_220_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hdc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_220_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_220_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hdd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_221_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_221_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hdd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_221_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_221_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hde == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_222_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_222_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hde == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_222_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_222_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hdf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_223_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_223_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hdf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_223_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_223_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_224_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_224_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_224_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_224_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_225_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_225_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_225_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_225_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_226_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_226_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_226_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_226_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_227_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_227_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_227_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_227_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_228_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_228_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_228_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_228_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_229_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_229_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_229_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_229_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_230_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_230_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_230_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_230_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_231_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_231_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_231_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_231_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_232_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_232_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_232_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_232_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_233_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_233_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'he9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_233_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_233_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hea == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_234_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_234_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hea == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_234_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_234_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'heb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_235_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_235_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'heb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_235_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_235_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hec == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_236_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_236_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hec == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_236_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_236_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hed == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_237_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_237_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hed == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_237_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_237_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hee == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_238_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_238_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hee == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_238_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_238_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hef == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_239_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_239_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hef == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_239_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_239_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_240_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_240_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_240_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_240_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_241_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_241_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_241_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_241_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_242_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_242_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_242_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_242_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_243_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_243_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_243_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_243_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_244_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_244_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_244_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_244_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_245_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_245_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_245_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_245_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_246_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_246_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_246_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_246_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_247_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_247_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_247_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_247_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_248_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_248_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_248_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_248_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_249_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_249_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hf9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_249_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_249_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfa == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_250_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_250_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfa == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_250_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_250_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_251_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_251_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_251_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_251_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_252_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_252_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_252_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_252_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_253_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_253_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_253_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_253_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfe == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_254_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_254_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hfe == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_254_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_254_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hff == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_255_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_255_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'hff == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_255_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_255_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h100 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_256_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_256_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h100 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_256_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_256_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h101 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_257_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_257_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h101 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_257_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_257_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h102 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_258_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_258_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h102 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_258_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_258_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h103 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_259_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_259_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h103 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_259_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_259_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h104 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_260_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_260_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h104 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_260_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_260_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h105 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_261_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_261_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h105 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_261_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_261_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h106 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_262_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_262_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h106 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_262_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_262_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h107 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_263_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_263_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h107 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_263_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_263_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h108 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_264_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_264_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h108 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_264_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_264_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h109 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_265_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_265_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h109 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_265_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_265_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_266_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_266_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_266_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_266_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_267_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_267_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_267_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_267_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_268_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_268_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_268_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_268_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_269_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_269_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_269_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_269_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_270_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_270_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_270_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_270_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_271_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_271_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h10f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_271_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_271_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h110 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_272_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_272_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h110 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_272_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_272_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h111 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_273_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_273_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h111 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_273_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_273_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h112 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_274_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_274_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h112 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_274_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_274_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h113 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_275_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_275_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h113 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_275_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_275_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h114 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_276_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_276_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h114 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_276_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_276_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h115 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_277_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_277_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h115 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_277_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_277_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h116 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_278_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_278_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h116 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_278_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_278_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h117 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_279_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_279_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h117 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_279_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_279_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h118 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_280_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_280_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h118 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_280_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_280_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h119 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_281_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_281_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h119 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_281_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_281_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_282_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_282_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_282_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_282_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_283_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_283_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_283_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_283_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_284_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_284_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_284_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_284_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_285_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_285_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_285_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_285_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_286_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_286_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_286_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_286_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_287_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_287_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h11f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_287_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_287_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h120 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_288_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_288_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h120 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_288_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_288_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h121 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_289_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_289_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h121 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_289_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_289_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h122 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_290_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_290_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h122 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_290_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_290_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h123 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_291_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_291_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h123 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_291_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_291_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h124 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_292_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_292_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h124 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_292_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_292_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h125 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_293_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_293_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h125 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_293_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_293_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h126 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_294_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_294_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h126 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_294_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_294_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h127 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_295_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_295_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h127 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_295_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_295_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h128 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_296_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_296_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h128 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_296_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_296_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h129 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_297_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_297_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h129 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_297_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_297_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_298_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_298_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_298_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_298_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_299_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_299_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_299_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_299_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_300_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_300_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_300_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_300_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_301_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_301_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_301_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_301_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_302_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_302_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_302_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_302_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_303_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_303_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h12f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_303_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_303_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h130 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_304_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_304_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h130 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_304_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_304_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h131 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_305_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_305_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h131 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_305_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_305_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h132 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_306_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_306_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h132 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_306_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_306_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h133 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_307_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_307_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h133 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_307_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_307_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h134 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_308_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_308_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h134 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_308_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_308_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h135 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_309_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_309_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h135 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_309_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_309_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h136 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_310_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_310_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h136 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_310_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_310_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h137 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_311_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_311_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h137 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_311_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_311_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h138 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_312_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_312_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h138 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_312_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_312_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h139 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_313_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_313_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h139 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_313_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_313_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_314_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_314_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_314_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_314_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_315_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_315_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_315_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_315_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_316_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_316_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_316_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_316_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_317_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_317_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_317_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_317_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_318_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_318_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_318_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_318_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_319_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_319_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h13f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_319_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_319_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h140 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_320_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_320_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h140 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_320_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_320_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h141 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_321_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_321_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h141 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_321_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_321_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h142 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_322_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_322_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h142 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_322_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_322_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h143 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_323_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_323_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h143 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_323_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_323_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h144 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_324_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_324_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h144 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_324_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_324_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h145 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_325_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_325_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h145 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_325_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_325_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h146 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_326_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_326_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h146 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_326_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_326_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h147 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_327_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_327_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h147 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_327_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_327_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h148 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_328_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_328_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h148 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_328_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_328_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h149 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_329_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_329_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h149 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_329_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_329_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_330_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_330_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_330_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_330_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_331_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_331_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_331_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_331_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_332_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_332_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_332_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_332_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_333_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_333_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_333_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_333_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_334_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_334_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_334_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_334_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_335_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_335_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h14f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_335_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_335_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h150 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_336_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_336_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h150 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_336_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_336_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h151 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_337_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_337_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h151 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_337_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_337_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h152 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_338_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_338_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h152 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_338_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_338_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h153 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_339_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_339_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h153 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_339_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_339_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h154 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_340_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_340_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h154 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_340_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_340_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h155 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_341_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_341_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h155 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_341_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_341_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h156 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_342_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_342_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h156 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_342_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_342_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h157 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_343_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_343_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h157 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_343_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_343_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h158 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_344_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_344_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h158 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_344_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_344_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h159 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_345_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_345_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h159 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_345_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_345_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_346_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_346_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_346_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_346_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_347_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_347_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_347_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_347_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_348_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_348_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_348_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_348_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_349_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_349_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_349_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_349_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_350_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_350_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_350_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_350_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_351_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_351_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h15f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_351_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_351_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h160 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_352_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_352_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h160 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_352_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_352_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h161 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_353_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_353_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h161 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_353_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_353_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h162 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_354_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_354_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h162 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_354_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_354_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h163 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_355_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_355_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h163 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_355_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_355_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h164 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_356_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_356_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h164 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_356_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_356_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h165 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_357_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_357_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h165 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_357_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_357_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h166 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_358_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_358_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h166 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_358_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_358_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h167 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_359_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_359_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h167 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_359_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_359_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h168 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_360_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_360_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h168 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_360_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_360_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h169 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_361_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_361_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h169 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_361_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_361_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_362_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_362_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_362_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_362_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_363_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_363_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_363_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_363_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_364_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_364_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_364_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_364_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_365_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_365_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_365_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_365_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_366_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_366_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_366_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_366_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_367_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_367_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h16f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_367_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_367_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h170 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_368_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_368_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h170 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_368_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_368_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h171 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_369_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_369_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h171 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_369_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_369_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h172 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_370_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_370_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h172 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_370_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_370_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h173 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_371_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_371_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h173 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_371_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_371_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h174 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_372_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_372_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h174 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_372_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_372_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h175 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_373_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_373_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h175 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_373_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_373_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h176 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_374_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_374_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h176 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_374_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_374_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h177 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_375_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_375_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h177 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_375_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_375_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h178 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_376_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_376_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h178 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_376_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_376_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h179 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_377_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_377_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h179 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_377_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_377_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_378_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_378_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_378_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_378_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_379_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_379_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_379_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_379_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_380_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_380_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_380_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_380_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_381_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_381_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_381_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_381_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_382_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_382_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_382_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_382_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_383_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_383_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h17f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_383_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_383_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h180 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_384_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_384_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h180 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_384_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_384_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h181 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_385_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_385_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h181 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_385_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_385_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h182 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_386_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_386_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h182 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_386_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_386_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h183 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_387_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_387_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h183 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_387_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_387_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h184 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_388_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_388_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h184 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_388_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_388_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h185 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_389_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_389_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h185 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_389_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_389_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h186 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_390_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_390_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h186 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_390_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_390_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h187 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_391_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_391_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h187 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_391_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_391_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h188 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_392_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_392_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h188 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_392_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_392_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h189 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_393_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_393_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h189 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_393_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_393_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_394_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_394_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_394_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_394_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_395_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_395_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_395_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_395_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_396_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_396_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_396_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_396_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_397_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_397_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_397_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_397_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_398_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_398_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_398_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_398_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_399_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_399_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h18f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_399_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_399_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h190 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_400_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_400_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h190 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_400_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_400_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h191 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_401_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_401_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h191 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_401_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_401_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h192 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_402_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_402_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h192 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_402_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_402_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h193 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_403_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_403_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h193 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_403_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_403_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h194 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_404_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_404_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h194 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_404_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_404_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h195 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_405_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_405_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h195 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_405_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_405_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h196 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_406_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_406_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h196 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_406_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_406_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h197 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_407_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_407_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h197 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_407_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_407_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h198 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_408_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_408_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h198 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_408_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_408_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h199 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_409_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_409_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h199 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_409_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_409_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_410_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_410_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_410_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_410_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_411_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_411_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_411_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_411_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_412_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_412_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_412_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_412_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_413_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_413_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_413_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_413_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_414_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_414_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_414_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_414_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_415_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_415_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h19f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_415_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_415_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_416_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_416_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_416_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_416_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_417_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_417_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_417_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_417_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_418_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_418_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_418_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_418_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_419_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_419_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_419_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_419_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_420_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_420_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_420_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_420_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_421_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_421_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_421_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_421_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_422_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_422_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_422_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_422_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_423_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_423_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_423_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_423_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_424_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_424_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_424_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_424_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_425_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_425_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1a9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_425_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_425_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1aa == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_426_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_426_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1aa == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_426_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_426_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ab == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_427_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_427_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ab == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_427_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_427_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ac == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_428_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_428_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ac == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_428_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_428_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ad == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_429_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_429_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ad == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_429_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_429_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ae == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_430_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_430_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ae == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_430_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_430_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1af == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_431_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_431_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1af == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_431_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_431_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_432_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_432_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_432_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_432_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_433_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_433_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_433_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_433_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_434_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_434_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_434_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_434_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_435_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_435_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_435_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_435_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_436_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_436_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_436_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_436_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_437_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_437_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_437_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_437_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_438_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_438_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_438_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_438_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_439_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_439_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_439_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_439_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_440_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_440_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_440_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_440_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_441_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_441_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1b9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_441_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_441_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ba == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_442_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_442_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ba == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_442_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_442_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1bb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_443_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_443_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1bb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_443_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_443_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1bc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_444_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_444_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1bc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_444_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_444_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1bd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_445_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_445_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1bd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_445_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_445_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1be == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_446_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_446_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1be == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_446_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_446_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1bf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_447_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_447_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1bf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_447_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_447_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_448_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_448_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_448_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_448_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_449_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_449_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_449_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_449_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_450_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_450_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_450_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_450_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_451_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_451_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_451_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_451_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_452_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_452_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_452_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_452_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_453_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_453_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_453_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_453_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_454_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_454_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_454_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_454_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_455_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_455_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_455_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_455_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_456_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_456_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_456_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_456_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_457_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_457_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1c9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_457_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_457_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ca == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_458_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_458_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ca == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_458_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_458_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1cb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_459_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_459_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1cb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_459_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_459_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1cc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_460_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_460_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1cc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_460_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_460_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1cd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_461_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_461_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1cd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_461_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_461_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ce == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_462_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_462_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ce == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_462_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_462_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1cf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_463_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_463_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1cf == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_463_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_463_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_464_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_464_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_464_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_464_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_465_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_465_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_465_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_465_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_466_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_466_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_466_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_466_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_467_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_467_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_467_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_467_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_468_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_468_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_468_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_468_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_469_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_469_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_469_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_469_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_470_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_470_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_470_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_470_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_471_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_471_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_471_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_471_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_472_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_472_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_472_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_472_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_473_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_473_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1d9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_473_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_473_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1da == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_474_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_474_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1da == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_474_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_474_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1db == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_475_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_475_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1db == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_475_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_475_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1dc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_476_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_476_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1dc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_476_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_476_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1dd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_477_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_477_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1dd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_477_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_477_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1de == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_478_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_478_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1de == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_478_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_478_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1df == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_479_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_479_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1df == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_479_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_479_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_480_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_480_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_480_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_480_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_481_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_481_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_481_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_481_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_482_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_482_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_482_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_482_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_483_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_483_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_483_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_483_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_484_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_484_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_484_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_484_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_485_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_485_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_485_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_485_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_486_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_486_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_486_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_486_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_487_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_487_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_487_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_487_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_488_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_488_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_488_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_488_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_489_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_489_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1e9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_489_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_489_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ea == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_490_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_490_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ea == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_490_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_490_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1eb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_491_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_491_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1eb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_491_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_491_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ec == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_492_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_492_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ec == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_492_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_492_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ed == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_493_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_493_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ed == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_493_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_493_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ee == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_494_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_494_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ee == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_494_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_494_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ef == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_495_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_495_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ef == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_495_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_495_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_496_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_496_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f0 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_496_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_496_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_497_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_497_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f1 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_497_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_497_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_498_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_498_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f2 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_498_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_498_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_499_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_499_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f3 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_499_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_499_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_500_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_500_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f4 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_500_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_500_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_501_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_501_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f5 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_501_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_501_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_502_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_502_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f6 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_502_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_502_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_503_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_503_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f7 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_503_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_503_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_504_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_504_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f8 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_504_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_504_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_505_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_505_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1f9 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_505_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_505_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fa == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_506_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_506_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fa == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_506_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_506_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_507_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_507_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fb == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_507_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_507_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_508_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_508_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fc == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_508_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_508_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_509_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_509_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fd == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_509_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_509_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fe == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_510_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_510_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1fe == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_510_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_510_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ff == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_511_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_511_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h1ff == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_511_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_511_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h200 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_512_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_512_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h200 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_512_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_512_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h201 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_513_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_513_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h201 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_513_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_513_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h202 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_514_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_514_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h202 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_514_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_514_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h203 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_515_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_515_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h203 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_515_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_515_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h204 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_516_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_516_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h204 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_516_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_516_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h205 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_517_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_517_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h205 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_517_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_517_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h206 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_518_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_518_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h206 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_518_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_518_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h207 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_519_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_519_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h207 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_519_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_519_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h208 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_520_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_520_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h208 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_520_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_520_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h209 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_521_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_521_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h209 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_521_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_521_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_522_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_522_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_522_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_522_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_523_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_523_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_523_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_523_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_524_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_524_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_524_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_524_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_525_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_525_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_525_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_525_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_526_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_526_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_526_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_526_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_527_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_527_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h20f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_527_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_527_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h210 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_528_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_528_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h210 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_528_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_528_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h211 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_529_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_529_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h211 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_529_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_529_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h212 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_530_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_530_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h212 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_530_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_530_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h213 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_531_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_531_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h213 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_531_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_531_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h214 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_532_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_532_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h214 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_532_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_532_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h215 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_533_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_533_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h215 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_533_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_533_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h216 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_534_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_534_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h216 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_534_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_534_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h217 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_535_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_535_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h217 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_535_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_535_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h218 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_536_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_536_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h218 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_536_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_536_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h219 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_537_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_537_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h219 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_537_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_537_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_538_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_538_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_538_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_538_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_539_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_539_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_539_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_539_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_540_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_540_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_540_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_540_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_541_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_541_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_541_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_541_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_542_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_542_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_542_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_542_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_543_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_543_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h21f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_543_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_543_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h220 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_544_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_544_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h220 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_544_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_544_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h221 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_545_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_545_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h221 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_545_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_545_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h222 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_546_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_546_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h222 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_546_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_546_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h223 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_547_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_547_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h223 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_547_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_547_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h224 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_548_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_548_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h224 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_548_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_548_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h225 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_549_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_549_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h225 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_549_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_549_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h226 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_550_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_550_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h226 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_550_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_550_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h227 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_551_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_551_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h227 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_551_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_551_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h228 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_552_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_552_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h228 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_552_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_552_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h229 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_553_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_553_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h229 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_553_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_553_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_554_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_554_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_554_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_554_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_555_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_555_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_555_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_555_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_556_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_556_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_556_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_556_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_557_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_557_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_557_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_557_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_558_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_558_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_558_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_558_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_559_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_559_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h22f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_559_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_559_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h230 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_560_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_560_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h230 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_560_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_560_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h231 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_561_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_561_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h231 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_561_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_561_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h232 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_562_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_562_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h232 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_562_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_562_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h233 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_563_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_563_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h233 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_563_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_563_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h234 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_564_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_564_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h234 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_564_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_564_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h235 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_565_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_565_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h235 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_565_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_565_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h236 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_566_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_566_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h236 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_566_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_566_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h237 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_567_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_567_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h237 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_567_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_567_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h238 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_568_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_568_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h238 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_568_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_568_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h239 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_569_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_569_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h239 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_569_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_569_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_570_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_570_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_570_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_570_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_571_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_571_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_571_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_571_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_572_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_572_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_572_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_572_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_573_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_573_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_573_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_573_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_574_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_574_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_574_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_574_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_575_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_575_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h23f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_575_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_575_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h240 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_576_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_576_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h240 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_576_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_576_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h241 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_577_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_577_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h241 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_577_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_577_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h242 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_578_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_578_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h242 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_578_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_578_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h243 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_579_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_579_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h243 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_579_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_579_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h244 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_580_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_580_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h244 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_580_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_580_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h245 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_581_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_581_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h245 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_581_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_581_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h246 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_582_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_582_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h246 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_582_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_582_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h247 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_583_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_583_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h247 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_583_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_583_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h248 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_584_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_584_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h248 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_584_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_584_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h249 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_585_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_585_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h249 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_585_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_585_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_586_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_586_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_586_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_586_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_587_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_587_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_587_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_587_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_588_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_588_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_588_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_588_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_589_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_589_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_589_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_589_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_590_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_590_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_590_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_590_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_591_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_591_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h24f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_591_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_591_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h250 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_592_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_592_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h250 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_592_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_592_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h251 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_593_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_593_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h251 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_593_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_593_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h252 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_594_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_594_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h252 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_594_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_594_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h253 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_595_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_595_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h253 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_595_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_595_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h254 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_596_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_596_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h254 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_596_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_596_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h255 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_597_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_597_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h255 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_597_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_597_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h256 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_598_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_598_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h256 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_598_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_598_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h257 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_599_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_599_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h257 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_599_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_599_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h258 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_600_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_600_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h258 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_600_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_600_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h259 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_601_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_601_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h259 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_601_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_601_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_602_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_602_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_602_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_602_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_603_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_603_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_603_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_603_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_604_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_604_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_604_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_604_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_605_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_605_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_605_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_605_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_606_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_606_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_606_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_606_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_607_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_607_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h25f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_607_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_607_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h260 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_608_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_608_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h260 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_608_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_608_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h261 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_609_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_609_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h261 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_609_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_609_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h262 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_610_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_610_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h262 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_610_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_610_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h263 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_611_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_611_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h263 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_611_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_611_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h264 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_612_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_612_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h264 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_612_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_612_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h265 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_613_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_613_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h265 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_613_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_613_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h266 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_614_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_614_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h266 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_614_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_614_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h267 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_615_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_615_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h267 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_615_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_615_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h268 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_616_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_616_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h268 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_616_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_616_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h269 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_617_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_617_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h269 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_617_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_617_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_618_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_618_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_618_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_618_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_619_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_619_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_619_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_619_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_620_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_620_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_620_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_620_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_621_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_621_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_621_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_621_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_622_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_622_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_622_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_622_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_623_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_623_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h26f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_623_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_623_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h270 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_624_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_624_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h270 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_624_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_624_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h271 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_625_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_625_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h271 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_625_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_625_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h272 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_626_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_626_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h272 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_626_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_626_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h273 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_627_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_627_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h273 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_627_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_627_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h274 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_628_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_628_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h274 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_628_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_628_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h275 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_629_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_629_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h275 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_629_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_629_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h276 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_630_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_630_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h276 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_630_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_630_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h277 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_631_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_631_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h277 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_631_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_631_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h278 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_632_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_632_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h278 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_632_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_632_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h279 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_633_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_633_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h279 == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_633_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_633_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_634_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_634_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27a == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_634_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_634_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_635_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_635_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27b == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_635_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_635_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_636_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_636_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27c == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_636_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_636_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_637_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_637_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27d == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_637_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_637_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_638_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_638_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27e == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_638_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_638_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_639_r <= last_px_r; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_639_r <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    if (10'h27f == io_x[9:0]) begin // @[EdgeDetect.scala 61:18]
      px_buffer_639_g <= last_px_g; // @[EdgeDetect.scala 61:18]
    end else begin
      px_buffer_639_g <= 8'h0; // @[EdgeDetect.scala 31:26]
    end
    last_px_r <= io_px_in_r; // @[EdgeDetect.scala 62:13]
    last_px_g <= io_px_in_g; // @[EdgeDetect.scala 62:13]
    if (io_x >= 11'h1) begin // @[EdgeDetect.scala 53:20]
      REG <= _T_62; // @[EdgeDetect.scala 54:13]
    end
    if (io_x >= 11'h1) begin // @[EdgeDetect.scala 53:20]
      REG_1 <= _T_80; // @[EdgeDetect.scala 56:13]
    end
    if (io_x >= 11'h1) begin // @[EdgeDetect.scala 53:20]
      REG_3 <= _T_70; // @[EdgeDetect.scala 55:13]
    end
    if (io_x >= 11'h1) begin // @[EdgeDetect.scala 53:20]
      REG_4 <= _T_88; // @[EdgeDetect.scala 57:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  px_buffer_0_r = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  px_buffer_0_g = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  px_buffer_1_r = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  px_buffer_1_g = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  px_buffer_2_r = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  px_buffer_2_g = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  px_buffer_3_r = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  px_buffer_3_g = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  px_buffer_4_r = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  px_buffer_4_g = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  px_buffer_5_r = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  px_buffer_5_g = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  px_buffer_6_r = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  px_buffer_6_g = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  px_buffer_7_r = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  px_buffer_7_g = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  px_buffer_8_r = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  px_buffer_8_g = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  px_buffer_9_r = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  px_buffer_9_g = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  px_buffer_10_r = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  px_buffer_10_g = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  px_buffer_11_r = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  px_buffer_11_g = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  px_buffer_12_r = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  px_buffer_12_g = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  px_buffer_13_r = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  px_buffer_13_g = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  px_buffer_14_r = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  px_buffer_14_g = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  px_buffer_15_r = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  px_buffer_15_g = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  px_buffer_16_r = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  px_buffer_16_g = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  px_buffer_17_r = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  px_buffer_17_g = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  px_buffer_18_r = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  px_buffer_18_g = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  px_buffer_19_r = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  px_buffer_19_g = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  px_buffer_20_r = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  px_buffer_20_g = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  px_buffer_21_r = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  px_buffer_21_g = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  px_buffer_22_r = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  px_buffer_22_g = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  px_buffer_23_r = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  px_buffer_23_g = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  px_buffer_24_r = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  px_buffer_24_g = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  px_buffer_25_r = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  px_buffer_25_g = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  px_buffer_26_r = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  px_buffer_26_g = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  px_buffer_27_r = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  px_buffer_27_g = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  px_buffer_28_r = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  px_buffer_28_g = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  px_buffer_29_r = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  px_buffer_29_g = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  px_buffer_30_r = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  px_buffer_30_g = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  px_buffer_31_r = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  px_buffer_31_g = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  px_buffer_32_r = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  px_buffer_32_g = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  px_buffer_33_r = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  px_buffer_33_g = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  px_buffer_34_r = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  px_buffer_34_g = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  px_buffer_35_r = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  px_buffer_35_g = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  px_buffer_36_r = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  px_buffer_36_g = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  px_buffer_37_r = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  px_buffer_37_g = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  px_buffer_38_r = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  px_buffer_38_g = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  px_buffer_39_r = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  px_buffer_39_g = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  px_buffer_40_r = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  px_buffer_40_g = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  px_buffer_41_r = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  px_buffer_41_g = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  px_buffer_42_r = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  px_buffer_42_g = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  px_buffer_43_r = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  px_buffer_43_g = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  px_buffer_44_r = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  px_buffer_44_g = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  px_buffer_45_r = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  px_buffer_45_g = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  px_buffer_46_r = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  px_buffer_46_g = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  px_buffer_47_r = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  px_buffer_47_g = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  px_buffer_48_r = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  px_buffer_48_g = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  px_buffer_49_r = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  px_buffer_49_g = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  px_buffer_50_r = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  px_buffer_50_g = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  px_buffer_51_r = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  px_buffer_51_g = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  px_buffer_52_r = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  px_buffer_52_g = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  px_buffer_53_r = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  px_buffer_53_g = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  px_buffer_54_r = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  px_buffer_54_g = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  px_buffer_55_r = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  px_buffer_55_g = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  px_buffer_56_r = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  px_buffer_56_g = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  px_buffer_57_r = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  px_buffer_57_g = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  px_buffer_58_r = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  px_buffer_58_g = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  px_buffer_59_r = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  px_buffer_59_g = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  px_buffer_60_r = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  px_buffer_60_g = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  px_buffer_61_r = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  px_buffer_61_g = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  px_buffer_62_r = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  px_buffer_62_g = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  px_buffer_63_r = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  px_buffer_63_g = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  px_buffer_64_r = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  px_buffer_64_g = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  px_buffer_65_r = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  px_buffer_65_g = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  px_buffer_66_r = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  px_buffer_66_g = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  px_buffer_67_r = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  px_buffer_67_g = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  px_buffer_68_r = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  px_buffer_68_g = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  px_buffer_69_r = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  px_buffer_69_g = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  px_buffer_70_r = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  px_buffer_70_g = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  px_buffer_71_r = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  px_buffer_71_g = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  px_buffer_72_r = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  px_buffer_72_g = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  px_buffer_73_r = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  px_buffer_73_g = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  px_buffer_74_r = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  px_buffer_74_g = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  px_buffer_75_r = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  px_buffer_75_g = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  px_buffer_76_r = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  px_buffer_76_g = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  px_buffer_77_r = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  px_buffer_77_g = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  px_buffer_78_r = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  px_buffer_78_g = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  px_buffer_79_r = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  px_buffer_79_g = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  px_buffer_80_r = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  px_buffer_80_g = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  px_buffer_81_r = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  px_buffer_81_g = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  px_buffer_82_r = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  px_buffer_82_g = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  px_buffer_83_r = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  px_buffer_83_g = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  px_buffer_84_r = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  px_buffer_84_g = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  px_buffer_85_r = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  px_buffer_85_g = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  px_buffer_86_r = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  px_buffer_86_g = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  px_buffer_87_r = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  px_buffer_87_g = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  px_buffer_88_r = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  px_buffer_88_g = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  px_buffer_89_r = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  px_buffer_89_g = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  px_buffer_90_r = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  px_buffer_90_g = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  px_buffer_91_r = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  px_buffer_91_g = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  px_buffer_92_r = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  px_buffer_92_g = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  px_buffer_93_r = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  px_buffer_93_g = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  px_buffer_94_r = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  px_buffer_94_g = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  px_buffer_95_r = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  px_buffer_95_g = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  px_buffer_96_r = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  px_buffer_96_g = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  px_buffer_97_r = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  px_buffer_97_g = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  px_buffer_98_r = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  px_buffer_98_g = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  px_buffer_99_r = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  px_buffer_99_g = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  px_buffer_100_r = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  px_buffer_100_g = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  px_buffer_101_r = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  px_buffer_101_g = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  px_buffer_102_r = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  px_buffer_102_g = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  px_buffer_103_r = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  px_buffer_103_g = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  px_buffer_104_r = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  px_buffer_104_g = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  px_buffer_105_r = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  px_buffer_105_g = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  px_buffer_106_r = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  px_buffer_106_g = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  px_buffer_107_r = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  px_buffer_107_g = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  px_buffer_108_r = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  px_buffer_108_g = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  px_buffer_109_r = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  px_buffer_109_g = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  px_buffer_110_r = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  px_buffer_110_g = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  px_buffer_111_r = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  px_buffer_111_g = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  px_buffer_112_r = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  px_buffer_112_g = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  px_buffer_113_r = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  px_buffer_113_g = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  px_buffer_114_r = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  px_buffer_114_g = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  px_buffer_115_r = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  px_buffer_115_g = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  px_buffer_116_r = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  px_buffer_116_g = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  px_buffer_117_r = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  px_buffer_117_g = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  px_buffer_118_r = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  px_buffer_118_g = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  px_buffer_119_r = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  px_buffer_119_g = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  px_buffer_120_r = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  px_buffer_120_g = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  px_buffer_121_r = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  px_buffer_121_g = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  px_buffer_122_r = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  px_buffer_122_g = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  px_buffer_123_r = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  px_buffer_123_g = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  px_buffer_124_r = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  px_buffer_124_g = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  px_buffer_125_r = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  px_buffer_125_g = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  px_buffer_126_r = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  px_buffer_126_g = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  px_buffer_127_r = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  px_buffer_127_g = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  px_buffer_128_r = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  px_buffer_128_g = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  px_buffer_129_r = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  px_buffer_129_g = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  px_buffer_130_r = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  px_buffer_130_g = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  px_buffer_131_r = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  px_buffer_131_g = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  px_buffer_132_r = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  px_buffer_132_g = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  px_buffer_133_r = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  px_buffer_133_g = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  px_buffer_134_r = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  px_buffer_134_g = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  px_buffer_135_r = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  px_buffer_135_g = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  px_buffer_136_r = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  px_buffer_136_g = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  px_buffer_137_r = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  px_buffer_137_g = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  px_buffer_138_r = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  px_buffer_138_g = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  px_buffer_139_r = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  px_buffer_139_g = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  px_buffer_140_r = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  px_buffer_140_g = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  px_buffer_141_r = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  px_buffer_141_g = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  px_buffer_142_r = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  px_buffer_142_g = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  px_buffer_143_r = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  px_buffer_143_g = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  px_buffer_144_r = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  px_buffer_144_g = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  px_buffer_145_r = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  px_buffer_145_g = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  px_buffer_146_r = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  px_buffer_146_g = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  px_buffer_147_r = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  px_buffer_147_g = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  px_buffer_148_r = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  px_buffer_148_g = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  px_buffer_149_r = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  px_buffer_149_g = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  px_buffer_150_r = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  px_buffer_150_g = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  px_buffer_151_r = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  px_buffer_151_g = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  px_buffer_152_r = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  px_buffer_152_g = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  px_buffer_153_r = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  px_buffer_153_g = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  px_buffer_154_r = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  px_buffer_154_g = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  px_buffer_155_r = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  px_buffer_155_g = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  px_buffer_156_r = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  px_buffer_156_g = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  px_buffer_157_r = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  px_buffer_157_g = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  px_buffer_158_r = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  px_buffer_158_g = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  px_buffer_159_r = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  px_buffer_159_g = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  px_buffer_160_r = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  px_buffer_160_g = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  px_buffer_161_r = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  px_buffer_161_g = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  px_buffer_162_r = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  px_buffer_162_g = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  px_buffer_163_r = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  px_buffer_163_g = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  px_buffer_164_r = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  px_buffer_164_g = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  px_buffer_165_r = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  px_buffer_165_g = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  px_buffer_166_r = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  px_buffer_166_g = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  px_buffer_167_r = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  px_buffer_167_g = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  px_buffer_168_r = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  px_buffer_168_g = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  px_buffer_169_r = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  px_buffer_169_g = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  px_buffer_170_r = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  px_buffer_170_g = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  px_buffer_171_r = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  px_buffer_171_g = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  px_buffer_172_r = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  px_buffer_172_g = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  px_buffer_173_r = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  px_buffer_173_g = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  px_buffer_174_r = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  px_buffer_174_g = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  px_buffer_175_r = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  px_buffer_175_g = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  px_buffer_176_r = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  px_buffer_176_g = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  px_buffer_177_r = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  px_buffer_177_g = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  px_buffer_178_r = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  px_buffer_178_g = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  px_buffer_179_r = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  px_buffer_179_g = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  px_buffer_180_r = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  px_buffer_180_g = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  px_buffer_181_r = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  px_buffer_181_g = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  px_buffer_182_r = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  px_buffer_182_g = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  px_buffer_183_r = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  px_buffer_183_g = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  px_buffer_184_r = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  px_buffer_184_g = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  px_buffer_185_r = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  px_buffer_185_g = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  px_buffer_186_r = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  px_buffer_186_g = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  px_buffer_187_r = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  px_buffer_187_g = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  px_buffer_188_r = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  px_buffer_188_g = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  px_buffer_189_r = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  px_buffer_189_g = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  px_buffer_190_r = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  px_buffer_190_g = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  px_buffer_191_r = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  px_buffer_191_g = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  px_buffer_192_r = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  px_buffer_192_g = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  px_buffer_193_r = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  px_buffer_193_g = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  px_buffer_194_r = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  px_buffer_194_g = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  px_buffer_195_r = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  px_buffer_195_g = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  px_buffer_196_r = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  px_buffer_196_g = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  px_buffer_197_r = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  px_buffer_197_g = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  px_buffer_198_r = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  px_buffer_198_g = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  px_buffer_199_r = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  px_buffer_199_g = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  px_buffer_200_r = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  px_buffer_200_g = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  px_buffer_201_r = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  px_buffer_201_g = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  px_buffer_202_r = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  px_buffer_202_g = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  px_buffer_203_r = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  px_buffer_203_g = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  px_buffer_204_r = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  px_buffer_204_g = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  px_buffer_205_r = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  px_buffer_205_g = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  px_buffer_206_r = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  px_buffer_206_g = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  px_buffer_207_r = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  px_buffer_207_g = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  px_buffer_208_r = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  px_buffer_208_g = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  px_buffer_209_r = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  px_buffer_209_g = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  px_buffer_210_r = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  px_buffer_210_g = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  px_buffer_211_r = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  px_buffer_211_g = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  px_buffer_212_r = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  px_buffer_212_g = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  px_buffer_213_r = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  px_buffer_213_g = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  px_buffer_214_r = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  px_buffer_214_g = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  px_buffer_215_r = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  px_buffer_215_g = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  px_buffer_216_r = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  px_buffer_216_g = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  px_buffer_217_r = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  px_buffer_217_g = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  px_buffer_218_r = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  px_buffer_218_g = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  px_buffer_219_r = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  px_buffer_219_g = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  px_buffer_220_r = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  px_buffer_220_g = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  px_buffer_221_r = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  px_buffer_221_g = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  px_buffer_222_r = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  px_buffer_222_g = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  px_buffer_223_r = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  px_buffer_223_g = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  px_buffer_224_r = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  px_buffer_224_g = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  px_buffer_225_r = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  px_buffer_225_g = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  px_buffer_226_r = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  px_buffer_226_g = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  px_buffer_227_r = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  px_buffer_227_g = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  px_buffer_228_r = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  px_buffer_228_g = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  px_buffer_229_r = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  px_buffer_229_g = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  px_buffer_230_r = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  px_buffer_230_g = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  px_buffer_231_r = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  px_buffer_231_g = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  px_buffer_232_r = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  px_buffer_232_g = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  px_buffer_233_r = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  px_buffer_233_g = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  px_buffer_234_r = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  px_buffer_234_g = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  px_buffer_235_r = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  px_buffer_235_g = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  px_buffer_236_r = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  px_buffer_236_g = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  px_buffer_237_r = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  px_buffer_237_g = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  px_buffer_238_r = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  px_buffer_238_g = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  px_buffer_239_r = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  px_buffer_239_g = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  px_buffer_240_r = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  px_buffer_240_g = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  px_buffer_241_r = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  px_buffer_241_g = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  px_buffer_242_r = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  px_buffer_242_g = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  px_buffer_243_r = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  px_buffer_243_g = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  px_buffer_244_r = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  px_buffer_244_g = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  px_buffer_245_r = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  px_buffer_245_g = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  px_buffer_246_r = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  px_buffer_246_g = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  px_buffer_247_r = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  px_buffer_247_g = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  px_buffer_248_r = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  px_buffer_248_g = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  px_buffer_249_r = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  px_buffer_249_g = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  px_buffer_250_r = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  px_buffer_250_g = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  px_buffer_251_r = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  px_buffer_251_g = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  px_buffer_252_r = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  px_buffer_252_g = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  px_buffer_253_r = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  px_buffer_253_g = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  px_buffer_254_r = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  px_buffer_254_g = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  px_buffer_255_r = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  px_buffer_255_g = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  px_buffer_256_r = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  px_buffer_256_g = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  px_buffer_257_r = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  px_buffer_257_g = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  px_buffer_258_r = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  px_buffer_258_g = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  px_buffer_259_r = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  px_buffer_259_g = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  px_buffer_260_r = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  px_buffer_260_g = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  px_buffer_261_r = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  px_buffer_261_g = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  px_buffer_262_r = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  px_buffer_262_g = _RAND_525[7:0];
  _RAND_526 = {1{`RANDOM}};
  px_buffer_263_r = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  px_buffer_263_g = _RAND_527[7:0];
  _RAND_528 = {1{`RANDOM}};
  px_buffer_264_r = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  px_buffer_264_g = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  px_buffer_265_r = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  px_buffer_265_g = _RAND_531[7:0];
  _RAND_532 = {1{`RANDOM}};
  px_buffer_266_r = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  px_buffer_266_g = _RAND_533[7:0];
  _RAND_534 = {1{`RANDOM}};
  px_buffer_267_r = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  px_buffer_267_g = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  px_buffer_268_r = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  px_buffer_268_g = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  px_buffer_269_r = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  px_buffer_269_g = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  px_buffer_270_r = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  px_buffer_270_g = _RAND_541[7:0];
  _RAND_542 = {1{`RANDOM}};
  px_buffer_271_r = _RAND_542[7:0];
  _RAND_543 = {1{`RANDOM}};
  px_buffer_271_g = _RAND_543[7:0];
  _RAND_544 = {1{`RANDOM}};
  px_buffer_272_r = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  px_buffer_272_g = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  px_buffer_273_r = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  px_buffer_273_g = _RAND_547[7:0];
  _RAND_548 = {1{`RANDOM}};
  px_buffer_274_r = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  px_buffer_274_g = _RAND_549[7:0];
  _RAND_550 = {1{`RANDOM}};
  px_buffer_275_r = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  px_buffer_275_g = _RAND_551[7:0];
  _RAND_552 = {1{`RANDOM}};
  px_buffer_276_r = _RAND_552[7:0];
  _RAND_553 = {1{`RANDOM}};
  px_buffer_276_g = _RAND_553[7:0];
  _RAND_554 = {1{`RANDOM}};
  px_buffer_277_r = _RAND_554[7:0];
  _RAND_555 = {1{`RANDOM}};
  px_buffer_277_g = _RAND_555[7:0];
  _RAND_556 = {1{`RANDOM}};
  px_buffer_278_r = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  px_buffer_278_g = _RAND_557[7:0];
  _RAND_558 = {1{`RANDOM}};
  px_buffer_279_r = _RAND_558[7:0];
  _RAND_559 = {1{`RANDOM}};
  px_buffer_279_g = _RAND_559[7:0];
  _RAND_560 = {1{`RANDOM}};
  px_buffer_280_r = _RAND_560[7:0];
  _RAND_561 = {1{`RANDOM}};
  px_buffer_280_g = _RAND_561[7:0];
  _RAND_562 = {1{`RANDOM}};
  px_buffer_281_r = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  px_buffer_281_g = _RAND_563[7:0];
  _RAND_564 = {1{`RANDOM}};
  px_buffer_282_r = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  px_buffer_282_g = _RAND_565[7:0];
  _RAND_566 = {1{`RANDOM}};
  px_buffer_283_r = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  px_buffer_283_g = _RAND_567[7:0];
  _RAND_568 = {1{`RANDOM}};
  px_buffer_284_r = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  px_buffer_284_g = _RAND_569[7:0];
  _RAND_570 = {1{`RANDOM}};
  px_buffer_285_r = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  px_buffer_285_g = _RAND_571[7:0];
  _RAND_572 = {1{`RANDOM}};
  px_buffer_286_r = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  px_buffer_286_g = _RAND_573[7:0];
  _RAND_574 = {1{`RANDOM}};
  px_buffer_287_r = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  px_buffer_287_g = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  px_buffer_288_r = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  px_buffer_288_g = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  px_buffer_289_r = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  px_buffer_289_g = _RAND_579[7:0];
  _RAND_580 = {1{`RANDOM}};
  px_buffer_290_r = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  px_buffer_290_g = _RAND_581[7:0];
  _RAND_582 = {1{`RANDOM}};
  px_buffer_291_r = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  px_buffer_291_g = _RAND_583[7:0];
  _RAND_584 = {1{`RANDOM}};
  px_buffer_292_r = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  px_buffer_292_g = _RAND_585[7:0];
  _RAND_586 = {1{`RANDOM}};
  px_buffer_293_r = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  px_buffer_293_g = _RAND_587[7:0];
  _RAND_588 = {1{`RANDOM}};
  px_buffer_294_r = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  px_buffer_294_g = _RAND_589[7:0];
  _RAND_590 = {1{`RANDOM}};
  px_buffer_295_r = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  px_buffer_295_g = _RAND_591[7:0];
  _RAND_592 = {1{`RANDOM}};
  px_buffer_296_r = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  px_buffer_296_g = _RAND_593[7:0];
  _RAND_594 = {1{`RANDOM}};
  px_buffer_297_r = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  px_buffer_297_g = _RAND_595[7:0];
  _RAND_596 = {1{`RANDOM}};
  px_buffer_298_r = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  px_buffer_298_g = _RAND_597[7:0];
  _RAND_598 = {1{`RANDOM}};
  px_buffer_299_r = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  px_buffer_299_g = _RAND_599[7:0];
  _RAND_600 = {1{`RANDOM}};
  px_buffer_300_r = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  px_buffer_300_g = _RAND_601[7:0];
  _RAND_602 = {1{`RANDOM}};
  px_buffer_301_r = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  px_buffer_301_g = _RAND_603[7:0];
  _RAND_604 = {1{`RANDOM}};
  px_buffer_302_r = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  px_buffer_302_g = _RAND_605[7:0];
  _RAND_606 = {1{`RANDOM}};
  px_buffer_303_r = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  px_buffer_303_g = _RAND_607[7:0];
  _RAND_608 = {1{`RANDOM}};
  px_buffer_304_r = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  px_buffer_304_g = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  px_buffer_305_r = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  px_buffer_305_g = _RAND_611[7:0];
  _RAND_612 = {1{`RANDOM}};
  px_buffer_306_r = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  px_buffer_306_g = _RAND_613[7:0];
  _RAND_614 = {1{`RANDOM}};
  px_buffer_307_r = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  px_buffer_307_g = _RAND_615[7:0];
  _RAND_616 = {1{`RANDOM}};
  px_buffer_308_r = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  px_buffer_308_g = _RAND_617[7:0];
  _RAND_618 = {1{`RANDOM}};
  px_buffer_309_r = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  px_buffer_309_g = _RAND_619[7:0];
  _RAND_620 = {1{`RANDOM}};
  px_buffer_310_r = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  px_buffer_310_g = _RAND_621[7:0];
  _RAND_622 = {1{`RANDOM}};
  px_buffer_311_r = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  px_buffer_311_g = _RAND_623[7:0];
  _RAND_624 = {1{`RANDOM}};
  px_buffer_312_r = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  px_buffer_312_g = _RAND_625[7:0];
  _RAND_626 = {1{`RANDOM}};
  px_buffer_313_r = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  px_buffer_313_g = _RAND_627[7:0];
  _RAND_628 = {1{`RANDOM}};
  px_buffer_314_r = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  px_buffer_314_g = _RAND_629[7:0];
  _RAND_630 = {1{`RANDOM}};
  px_buffer_315_r = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  px_buffer_315_g = _RAND_631[7:0];
  _RAND_632 = {1{`RANDOM}};
  px_buffer_316_r = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  px_buffer_316_g = _RAND_633[7:0];
  _RAND_634 = {1{`RANDOM}};
  px_buffer_317_r = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  px_buffer_317_g = _RAND_635[7:0];
  _RAND_636 = {1{`RANDOM}};
  px_buffer_318_r = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  px_buffer_318_g = _RAND_637[7:0];
  _RAND_638 = {1{`RANDOM}};
  px_buffer_319_r = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  px_buffer_319_g = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  px_buffer_320_r = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  px_buffer_320_g = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  px_buffer_321_r = _RAND_642[7:0];
  _RAND_643 = {1{`RANDOM}};
  px_buffer_321_g = _RAND_643[7:0];
  _RAND_644 = {1{`RANDOM}};
  px_buffer_322_r = _RAND_644[7:0];
  _RAND_645 = {1{`RANDOM}};
  px_buffer_322_g = _RAND_645[7:0];
  _RAND_646 = {1{`RANDOM}};
  px_buffer_323_r = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  px_buffer_323_g = _RAND_647[7:0];
  _RAND_648 = {1{`RANDOM}};
  px_buffer_324_r = _RAND_648[7:0];
  _RAND_649 = {1{`RANDOM}};
  px_buffer_324_g = _RAND_649[7:0];
  _RAND_650 = {1{`RANDOM}};
  px_buffer_325_r = _RAND_650[7:0];
  _RAND_651 = {1{`RANDOM}};
  px_buffer_325_g = _RAND_651[7:0];
  _RAND_652 = {1{`RANDOM}};
  px_buffer_326_r = _RAND_652[7:0];
  _RAND_653 = {1{`RANDOM}};
  px_buffer_326_g = _RAND_653[7:0];
  _RAND_654 = {1{`RANDOM}};
  px_buffer_327_r = _RAND_654[7:0];
  _RAND_655 = {1{`RANDOM}};
  px_buffer_327_g = _RAND_655[7:0];
  _RAND_656 = {1{`RANDOM}};
  px_buffer_328_r = _RAND_656[7:0];
  _RAND_657 = {1{`RANDOM}};
  px_buffer_328_g = _RAND_657[7:0];
  _RAND_658 = {1{`RANDOM}};
  px_buffer_329_r = _RAND_658[7:0];
  _RAND_659 = {1{`RANDOM}};
  px_buffer_329_g = _RAND_659[7:0];
  _RAND_660 = {1{`RANDOM}};
  px_buffer_330_r = _RAND_660[7:0];
  _RAND_661 = {1{`RANDOM}};
  px_buffer_330_g = _RAND_661[7:0];
  _RAND_662 = {1{`RANDOM}};
  px_buffer_331_r = _RAND_662[7:0];
  _RAND_663 = {1{`RANDOM}};
  px_buffer_331_g = _RAND_663[7:0];
  _RAND_664 = {1{`RANDOM}};
  px_buffer_332_r = _RAND_664[7:0];
  _RAND_665 = {1{`RANDOM}};
  px_buffer_332_g = _RAND_665[7:0];
  _RAND_666 = {1{`RANDOM}};
  px_buffer_333_r = _RAND_666[7:0];
  _RAND_667 = {1{`RANDOM}};
  px_buffer_333_g = _RAND_667[7:0];
  _RAND_668 = {1{`RANDOM}};
  px_buffer_334_r = _RAND_668[7:0];
  _RAND_669 = {1{`RANDOM}};
  px_buffer_334_g = _RAND_669[7:0];
  _RAND_670 = {1{`RANDOM}};
  px_buffer_335_r = _RAND_670[7:0];
  _RAND_671 = {1{`RANDOM}};
  px_buffer_335_g = _RAND_671[7:0];
  _RAND_672 = {1{`RANDOM}};
  px_buffer_336_r = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  px_buffer_336_g = _RAND_673[7:0];
  _RAND_674 = {1{`RANDOM}};
  px_buffer_337_r = _RAND_674[7:0];
  _RAND_675 = {1{`RANDOM}};
  px_buffer_337_g = _RAND_675[7:0];
  _RAND_676 = {1{`RANDOM}};
  px_buffer_338_r = _RAND_676[7:0];
  _RAND_677 = {1{`RANDOM}};
  px_buffer_338_g = _RAND_677[7:0];
  _RAND_678 = {1{`RANDOM}};
  px_buffer_339_r = _RAND_678[7:0];
  _RAND_679 = {1{`RANDOM}};
  px_buffer_339_g = _RAND_679[7:0];
  _RAND_680 = {1{`RANDOM}};
  px_buffer_340_r = _RAND_680[7:0];
  _RAND_681 = {1{`RANDOM}};
  px_buffer_340_g = _RAND_681[7:0];
  _RAND_682 = {1{`RANDOM}};
  px_buffer_341_r = _RAND_682[7:0];
  _RAND_683 = {1{`RANDOM}};
  px_buffer_341_g = _RAND_683[7:0];
  _RAND_684 = {1{`RANDOM}};
  px_buffer_342_r = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  px_buffer_342_g = _RAND_685[7:0];
  _RAND_686 = {1{`RANDOM}};
  px_buffer_343_r = _RAND_686[7:0];
  _RAND_687 = {1{`RANDOM}};
  px_buffer_343_g = _RAND_687[7:0];
  _RAND_688 = {1{`RANDOM}};
  px_buffer_344_r = _RAND_688[7:0];
  _RAND_689 = {1{`RANDOM}};
  px_buffer_344_g = _RAND_689[7:0];
  _RAND_690 = {1{`RANDOM}};
  px_buffer_345_r = _RAND_690[7:0];
  _RAND_691 = {1{`RANDOM}};
  px_buffer_345_g = _RAND_691[7:0];
  _RAND_692 = {1{`RANDOM}};
  px_buffer_346_r = _RAND_692[7:0];
  _RAND_693 = {1{`RANDOM}};
  px_buffer_346_g = _RAND_693[7:0];
  _RAND_694 = {1{`RANDOM}};
  px_buffer_347_r = _RAND_694[7:0];
  _RAND_695 = {1{`RANDOM}};
  px_buffer_347_g = _RAND_695[7:0];
  _RAND_696 = {1{`RANDOM}};
  px_buffer_348_r = _RAND_696[7:0];
  _RAND_697 = {1{`RANDOM}};
  px_buffer_348_g = _RAND_697[7:0];
  _RAND_698 = {1{`RANDOM}};
  px_buffer_349_r = _RAND_698[7:0];
  _RAND_699 = {1{`RANDOM}};
  px_buffer_349_g = _RAND_699[7:0];
  _RAND_700 = {1{`RANDOM}};
  px_buffer_350_r = _RAND_700[7:0];
  _RAND_701 = {1{`RANDOM}};
  px_buffer_350_g = _RAND_701[7:0];
  _RAND_702 = {1{`RANDOM}};
  px_buffer_351_r = _RAND_702[7:0];
  _RAND_703 = {1{`RANDOM}};
  px_buffer_351_g = _RAND_703[7:0];
  _RAND_704 = {1{`RANDOM}};
  px_buffer_352_r = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  px_buffer_352_g = _RAND_705[7:0];
  _RAND_706 = {1{`RANDOM}};
  px_buffer_353_r = _RAND_706[7:0];
  _RAND_707 = {1{`RANDOM}};
  px_buffer_353_g = _RAND_707[7:0];
  _RAND_708 = {1{`RANDOM}};
  px_buffer_354_r = _RAND_708[7:0];
  _RAND_709 = {1{`RANDOM}};
  px_buffer_354_g = _RAND_709[7:0];
  _RAND_710 = {1{`RANDOM}};
  px_buffer_355_r = _RAND_710[7:0];
  _RAND_711 = {1{`RANDOM}};
  px_buffer_355_g = _RAND_711[7:0];
  _RAND_712 = {1{`RANDOM}};
  px_buffer_356_r = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  px_buffer_356_g = _RAND_713[7:0];
  _RAND_714 = {1{`RANDOM}};
  px_buffer_357_r = _RAND_714[7:0];
  _RAND_715 = {1{`RANDOM}};
  px_buffer_357_g = _RAND_715[7:0];
  _RAND_716 = {1{`RANDOM}};
  px_buffer_358_r = _RAND_716[7:0];
  _RAND_717 = {1{`RANDOM}};
  px_buffer_358_g = _RAND_717[7:0];
  _RAND_718 = {1{`RANDOM}};
  px_buffer_359_r = _RAND_718[7:0];
  _RAND_719 = {1{`RANDOM}};
  px_buffer_359_g = _RAND_719[7:0];
  _RAND_720 = {1{`RANDOM}};
  px_buffer_360_r = _RAND_720[7:0];
  _RAND_721 = {1{`RANDOM}};
  px_buffer_360_g = _RAND_721[7:0];
  _RAND_722 = {1{`RANDOM}};
  px_buffer_361_r = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  px_buffer_361_g = _RAND_723[7:0];
  _RAND_724 = {1{`RANDOM}};
  px_buffer_362_r = _RAND_724[7:0];
  _RAND_725 = {1{`RANDOM}};
  px_buffer_362_g = _RAND_725[7:0];
  _RAND_726 = {1{`RANDOM}};
  px_buffer_363_r = _RAND_726[7:0];
  _RAND_727 = {1{`RANDOM}};
  px_buffer_363_g = _RAND_727[7:0];
  _RAND_728 = {1{`RANDOM}};
  px_buffer_364_r = _RAND_728[7:0];
  _RAND_729 = {1{`RANDOM}};
  px_buffer_364_g = _RAND_729[7:0];
  _RAND_730 = {1{`RANDOM}};
  px_buffer_365_r = _RAND_730[7:0];
  _RAND_731 = {1{`RANDOM}};
  px_buffer_365_g = _RAND_731[7:0];
  _RAND_732 = {1{`RANDOM}};
  px_buffer_366_r = _RAND_732[7:0];
  _RAND_733 = {1{`RANDOM}};
  px_buffer_366_g = _RAND_733[7:0];
  _RAND_734 = {1{`RANDOM}};
  px_buffer_367_r = _RAND_734[7:0];
  _RAND_735 = {1{`RANDOM}};
  px_buffer_367_g = _RAND_735[7:0];
  _RAND_736 = {1{`RANDOM}};
  px_buffer_368_r = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  px_buffer_368_g = _RAND_737[7:0];
  _RAND_738 = {1{`RANDOM}};
  px_buffer_369_r = _RAND_738[7:0];
  _RAND_739 = {1{`RANDOM}};
  px_buffer_369_g = _RAND_739[7:0];
  _RAND_740 = {1{`RANDOM}};
  px_buffer_370_r = _RAND_740[7:0];
  _RAND_741 = {1{`RANDOM}};
  px_buffer_370_g = _RAND_741[7:0];
  _RAND_742 = {1{`RANDOM}};
  px_buffer_371_r = _RAND_742[7:0];
  _RAND_743 = {1{`RANDOM}};
  px_buffer_371_g = _RAND_743[7:0];
  _RAND_744 = {1{`RANDOM}};
  px_buffer_372_r = _RAND_744[7:0];
  _RAND_745 = {1{`RANDOM}};
  px_buffer_372_g = _RAND_745[7:0];
  _RAND_746 = {1{`RANDOM}};
  px_buffer_373_r = _RAND_746[7:0];
  _RAND_747 = {1{`RANDOM}};
  px_buffer_373_g = _RAND_747[7:0];
  _RAND_748 = {1{`RANDOM}};
  px_buffer_374_r = _RAND_748[7:0];
  _RAND_749 = {1{`RANDOM}};
  px_buffer_374_g = _RAND_749[7:0];
  _RAND_750 = {1{`RANDOM}};
  px_buffer_375_r = _RAND_750[7:0];
  _RAND_751 = {1{`RANDOM}};
  px_buffer_375_g = _RAND_751[7:0];
  _RAND_752 = {1{`RANDOM}};
  px_buffer_376_r = _RAND_752[7:0];
  _RAND_753 = {1{`RANDOM}};
  px_buffer_376_g = _RAND_753[7:0];
  _RAND_754 = {1{`RANDOM}};
  px_buffer_377_r = _RAND_754[7:0];
  _RAND_755 = {1{`RANDOM}};
  px_buffer_377_g = _RAND_755[7:0];
  _RAND_756 = {1{`RANDOM}};
  px_buffer_378_r = _RAND_756[7:0];
  _RAND_757 = {1{`RANDOM}};
  px_buffer_378_g = _RAND_757[7:0];
  _RAND_758 = {1{`RANDOM}};
  px_buffer_379_r = _RAND_758[7:0];
  _RAND_759 = {1{`RANDOM}};
  px_buffer_379_g = _RAND_759[7:0];
  _RAND_760 = {1{`RANDOM}};
  px_buffer_380_r = _RAND_760[7:0];
  _RAND_761 = {1{`RANDOM}};
  px_buffer_380_g = _RAND_761[7:0];
  _RAND_762 = {1{`RANDOM}};
  px_buffer_381_r = _RAND_762[7:0];
  _RAND_763 = {1{`RANDOM}};
  px_buffer_381_g = _RAND_763[7:0];
  _RAND_764 = {1{`RANDOM}};
  px_buffer_382_r = _RAND_764[7:0];
  _RAND_765 = {1{`RANDOM}};
  px_buffer_382_g = _RAND_765[7:0];
  _RAND_766 = {1{`RANDOM}};
  px_buffer_383_r = _RAND_766[7:0];
  _RAND_767 = {1{`RANDOM}};
  px_buffer_383_g = _RAND_767[7:0];
  _RAND_768 = {1{`RANDOM}};
  px_buffer_384_r = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  px_buffer_384_g = _RAND_769[7:0];
  _RAND_770 = {1{`RANDOM}};
  px_buffer_385_r = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  px_buffer_385_g = _RAND_771[7:0];
  _RAND_772 = {1{`RANDOM}};
  px_buffer_386_r = _RAND_772[7:0];
  _RAND_773 = {1{`RANDOM}};
  px_buffer_386_g = _RAND_773[7:0];
  _RAND_774 = {1{`RANDOM}};
  px_buffer_387_r = _RAND_774[7:0];
  _RAND_775 = {1{`RANDOM}};
  px_buffer_387_g = _RAND_775[7:0];
  _RAND_776 = {1{`RANDOM}};
  px_buffer_388_r = _RAND_776[7:0];
  _RAND_777 = {1{`RANDOM}};
  px_buffer_388_g = _RAND_777[7:0];
  _RAND_778 = {1{`RANDOM}};
  px_buffer_389_r = _RAND_778[7:0];
  _RAND_779 = {1{`RANDOM}};
  px_buffer_389_g = _RAND_779[7:0];
  _RAND_780 = {1{`RANDOM}};
  px_buffer_390_r = _RAND_780[7:0];
  _RAND_781 = {1{`RANDOM}};
  px_buffer_390_g = _RAND_781[7:0];
  _RAND_782 = {1{`RANDOM}};
  px_buffer_391_r = _RAND_782[7:0];
  _RAND_783 = {1{`RANDOM}};
  px_buffer_391_g = _RAND_783[7:0];
  _RAND_784 = {1{`RANDOM}};
  px_buffer_392_r = _RAND_784[7:0];
  _RAND_785 = {1{`RANDOM}};
  px_buffer_392_g = _RAND_785[7:0];
  _RAND_786 = {1{`RANDOM}};
  px_buffer_393_r = _RAND_786[7:0];
  _RAND_787 = {1{`RANDOM}};
  px_buffer_393_g = _RAND_787[7:0];
  _RAND_788 = {1{`RANDOM}};
  px_buffer_394_r = _RAND_788[7:0];
  _RAND_789 = {1{`RANDOM}};
  px_buffer_394_g = _RAND_789[7:0];
  _RAND_790 = {1{`RANDOM}};
  px_buffer_395_r = _RAND_790[7:0];
  _RAND_791 = {1{`RANDOM}};
  px_buffer_395_g = _RAND_791[7:0];
  _RAND_792 = {1{`RANDOM}};
  px_buffer_396_r = _RAND_792[7:0];
  _RAND_793 = {1{`RANDOM}};
  px_buffer_396_g = _RAND_793[7:0];
  _RAND_794 = {1{`RANDOM}};
  px_buffer_397_r = _RAND_794[7:0];
  _RAND_795 = {1{`RANDOM}};
  px_buffer_397_g = _RAND_795[7:0];
  _RAND_796 = {1{`RANDOM}};
  px_buffer_398_r = _RAND_796[7:0];
  _RAND_797 = {1{`RANDOM}};
  px_buffer_398_g = _RAND_797[7:0];
  _RAND_798 = {1{`RANDOM}};
  px_buffer_399_r = _RAND_798[7:0];
  _RAND_799 = {1{`RANDOM}};
  px_buffer_399_g = _RAND_799[7:0];
  _RAND_800 = {1{`RANDOM}};
  px_buffer_400_r = _RAND_800[7:0];
  _RAND_801 = {1{`RANDOM}};
  px_buffer_400_g = _RAND_801[7:0];
  _RAND_802 = {1{`RANDOM}};
  px_buffer_401_r = _RAND_802[7:0];
  _RAND_803 = {1{`RANDOM}};
  px_buffer_401_g = _RAND_803[7:0];
  _RAND_804 = {1{`RANDOM}};
  px_buffer_402_r = _RAND_804[7:0];
  _RAND_805 = {1{`RANDOM}};
  px_buffer_402_g = _RAND_805[7:0];
  _RAND_806 = {1{`RANDOM}};
  px_buffer_403_r = _RAND_806[7:0];
  _RAND_807 = {1{`RANDOM}};
  px_buffer_403_g = _RAND_807[7:0];
  _RAND_808 = {1{`RANDOM}};
  px_buffer_404_r = _RAND_808[7:0];
  _RAND_809 = {1{`RANDOM}};
  px_buffer_404_g = _RAND_809[7:0];
  _RAND_810 = {1{`RANDOM}};
  px_buffer_405_r = _RAND_810[7:0];
  _RAND_811 = {1{`RANDOM}};
  px_buffer_405_g = _RAND_811[7:0];
  _RAND_812 = {1{`RANDOM}};
  px_buffer_406_r = _RAND_812[7:0];
  _RAND_813 = {1{`RANDOM}};
  px_buffer_406_g = _RAND_813[7:0];
  _RAND_814 = {1{`RANDOM}};
  px_buffer_407_r = _RAND_814[7:0];
  _RAND_815 = {1{`RANDOM}};
  px_buffer_407_g = _RAND_815[7:0];
  _RAND_816 = {1{`RANDOM}};
  px_buffer_408_r = _RAND_816[7:0];
  _RAND_817 = {1{`RANDOM}};
  px_buffer_408_g = _RAND_817[7:0];
  _RAND_818 = {1{`RANDOM}};
  px_buffer_409_r = _RAND_818[7:0];
  _RAND_819 = {1{`RANDOM}};
  px_buffer_409_g = _RAND_819[7:0];
  _RAND_820 = {1{`RANDOM}};
  px_buffer_410_r = _RAND_820[7:0];
  _RAND_821 = {1{`RANDOM}};
  px_buffer_410_g = _RAND_821[7:0];
  _RAND_822 = {1{`RANDOM}};
  px_buffer_411_r = _RAND_822[7:0];
  _RAND_823 = {1{`RANDOM}};
  px_buffer_411_g = _RAND_823[7:0];
  _RAND_824 = {1{`RANDOM}};
  px_buffer_412_r = _RAND_824[7:0];
  _RAND_825 = {1{`RANDOM}};
  px_buffer_412_g = _RAND_825[7:0];
  _RAND_826 = {1{`RANDOM}};
  px_buffer_413_r = _RAND_826[7:0];
  _RAND_827 = {1{`RANDOM}};
  px_buffer_413_g = _RAND_827[7:0];
  _RAND_828 = {1{`RANDOM}};
  px_buffer_414_r = _RAND_828[7:0];
  _RAND_829 = {1{`RANDOM}};
  px_buffer_414_g = _RAND_829[7:0];
  _RAND_830 = {1{`RANDOM}};
  px_buffer_415_r = _RAND_830[7:0];
  _RAND_831 = {1{`RANDOM}};
  px_buffer_415_g = _RAND_831[7:0];
  _RAND_832 = {1{`RANDOM}};
  px_buffer_416_r = _RAND_832[7:0];
  _RAND_833 = {1{`RANDOM}};
  px_buffer_416_g = _RAND_833[7:0];
  _RAND_834 = {1{`RANDOM}};
  px_buffer_417_r = _RAND_834[7:0];
  _RAND_835 = {1{`RANDOM}};
  px_buffer_417_g = _RAND_835[7:0];
  _RAND_836 = {1{`RANDOM}};
  px_buffer_418_r = _RAND_836[7:0];
  _RAND_837 = {1{`RANDOM}};
  px_buffer_418_g = _RAND_837[7:0];
  _RAND_838 = {1{`RANDOM}};
  px_buffer_419_r = _RAND_838[7:0];
  _RAND_839 = {1{`RANDOM}};
  px_buffer_419_g = _RAND_839[7:0];
  _RAND_840 = {1{`RANDOM}};
  px_buffer_420_r = _RAND_840[7:0];
  _RAND_841 = {1{`RANDOM}};
  px_buffer_420_g = _RAND_841[7:0];
  _RAND_842 = {1{`RANDOM}};
  px_buffer_421_r = _RAND_842[7:0];
  _RAND_843 = {1{`RANDOM}};
  px_buffer_421_g = _RAND_843[7:0];
  _RAND_844 = {1{`RANDOM}};
  px_buffer_422_r = _RAND_844[7:0];
  _RAND_845 = {1{`RANDOM}};
  px_buffer_422_g = _RAND_845[7:0];
  _RAND_846 = {1{`RANDOM}};
  px_buffer_423_r = _RAND_846[7:0];
  _RAND_847 = {1{`RANDOM}};
  px_buffer_423_g = _RAND_847[7:0];
  _RAND_848 = {1{`RANDOM}};
  px_buffer_424_r = _RAND_848[7:0];
  _RAND_849 = {1{`RANDOM}};
  px_buffer_424_g = _RAND_849[7:0];
  _RAND_850 = {1{`RANDOM}};
  px_buffer_425_r = _RAND_850[7:0];
  _RAND_851 = {1{`RANDOM}};
  px_buffer_425_g = _RAND_851[7:0];
  _RAND_852 = {1{`RANDOM}};
  px_buffer_426_r = _RAND_852[7:0];
  _RAND_853 = {1{`RANDOM}};
  px_buffer_426_g = _RAND_853[7:0];
  _RAND_854 = {1{`RANDOM}};
  px_buffer_427_r = _RAND_854[7:0];
  _RAND_855 = {1{`RANDOM}};
  px_buffer_427_g = _RAND_855[7:0];
  _RAND_856 = {1{`RANDOM}};
  px_buffer_428_r = _RAND_856[7:0];
  _RAND_857 = {1{`RANDOM}};
  px_buffer_428_g = _RAND_857[7:0];
  _RAND_858 = {1{`RANDOM}};
  px_buffer_429_r = _RAND_858[7:0];
  _RAND_859 = {1{`RANDOM}};
  px_buffer_429_g = _RAND_859[7:0];
  _RAND_860 = {1{`RANDOM}};
  px_buffer_430_r = _RAND_860[7:0];
  _RAND_861 = {1{`RANDOM}};
  px_buffer_430_g = _RAND_861[7:0];
  _RAND_862 = {1{`RANDOM}};
  px_buffer_431_r = _RAND_862[7:0];
  _RAND_863 = {1{`RANDOM}};
  px_buffer_431_g = _RAND_863[7:0];
  _RAND_864 = {1{`RANDOM}};
  px_buffer_432_r = _RAND_864[7:0];
  _RAND_865 = {1{`RANDOM}};
  px_buffer_432_g = _RAND_865[7:0];
  _RAND_866 = {1{`RANDOM}};
  px_buffer_433_r = _RAND_866[7:0];
  _RAND_867 = {1{`RANDOM}};
  px_buffer_433_g = _RAND_867[7:0];
  _RAND_868 = {1{`RANDOM}};
  px_buffer_434_r = _RAND_868[7:0];
  _RAND_869 = {1{`RANDOM}};
  px_buffer_434_g = _RAND_869[7:0];
  _RAND_870 = {1{`RANDOM}};
  px_buffer_435_r = _RAND_870[7:0];
  _RAND_871 = {1{`RANDOM}};
  px_buffer_435_g = _RAND_871[7:0];
  _RAND_872 = {1{`RANDOM}};
  px_buffer_436_r = _RAND_872[7:0];
  _RAND_873 = {1{`RANDOM}};
  px_buffer_436_g = _RAND_873[7:0];
  _RAND_874 = {1{`RANDOM}};
  px_buffer_437_r = _RAND_874[7:0];
  _RAND_875 = {1{`RANDOM}};
  px_buffer_437_g = _RAND_875[7:0];
  _RAND_876 = {1{`RANDOM}};
  px_buffer_438_r = _RAND_876[7:0];
  _RAND_877 = {1{`RANDOM}};
  px_buffer_438_g = _RAND_877[7:0];
  _RAND_878 = {1{`RANDOM}};
  px_buffer_439_r = _RAND_878[7:0];
  _RAND_879 = {1{`RANDOM}};
  px_buffer_439_g = _RAND_879[7:0];
  _RAND_880 = {1{`RANDOM}};
  px_buffer_440_r = _RAND_880[7:0];
  _RAND_881 = {1{`RANDOM}};
  px_buffer_440_g = _RAND_881[7:0];
  _RAND_882 = {1{`RANDOM}};
  px_buffer_441_r = _RAND_882[7:0];
  _RAND_883 = {1{`RANDOM}};
  px_buffer_441_g = _RAND_883[7:0];
  _RAND_884 = {1{`RANDOM}};
  px_buffer_442_r = _RAND_884[7:0];
  _RAND_885 = {1{`RANDOM}};
  px_buffer_442_g = _RAND_885[7:0];
  _RAND_886 = {1{`RANDOM}};
  px_buffer_443_r = _RAND_886[7:0];
  _RAND_887 = {1{`RANDOM}};
  px_buffer_443_g = _RAND_887[7:0];
  _RAND_888 = {1{`RANDOM}};
  px_buffer_444_r = _RAND_888[7:0];
  _RAND_889 = {1{`RANDOM}};
  px_buffer_444_g = _RAND_889[7:0];
  _RAND_890 = {1{`RANDOM}};
  px_buffer_445_r = _RAND_890[7:0];
  _RAND_891 = {1{`RANDOM}};
  px_buffer_445_g = _RAND_891[7:0];
  _RAND_892 = {1{`RANDOM}};
  px_buffer_446_r = _RAND_892[7:0];
  _RAND_893 = {1{`RANDOM}};
  px_buffer_446_g = _RAND_893[7:0];
  _RAND_894 = {1{`RANDOM}};
  px_buffer_447_r = _RAND_894[7:0];
  _RAND_895 = {1{`RANDOM}};
  px_buffer_447_g = _RAND_895[7:0];
  _RAND_896 = {1{`RANDOM}};
  px_buffer_448_r = _RAND_896[7:0];
  _RAND_897 = {1{`RANDOM}};
  px_buffer_448_g = _RAND_897[7:0];
  _RAND_898 = {1{`RANDOM}};
  px_buffer_449_r = _RAND_898[7:0];
  _RAND_899 = {1{`RANDOM}};
  px_buffer_449_g = _RAND_899[7:0];
  _RAND_900 = {1{`RANDOM}};
  px_buffer_450_r = _RAND_900[7:0];
  _RAND_901 = {1{`RANDOM}};
  px_buffer_450_g = _RAND_901[7:0];
  _RAND_902 = {1{`RANDOM}};
  px_buffer_451_r = _RAND_902[7:0];
  _RAND_903 = {1{`RANDOM}};
  px_buffer_451_g = _RAND_903[7:0];
  _RAND_904 = {1{`RANDOM}};
  px_buffer_452_r = _RAND_904[7:0];
  _RAND_905 = {1{`RANDOM}};
  px_buffer_452_g = _RAND_905[7:0];
  _RAND_906 = {1{`RANDOM}};
  px_buffer_453_r = _RAND_906[7:0];
  _RAND_907 = {1{`RANDOM}};
  px_buffer_453_g = _RAND_907[7:0];
  _RAND_908 = {1{`RANDOM}};
  px_buffer_454_r = _RAND_908[7:0];
  _RAND_909 = {1{`RANDOM}};
  px_buffer_454_g = _RAND_909[7:0];
  _RAND_910 = {1{`RANDOM}};
  px_buffer_455_r = _RAND_910[7:0];
  _RAND_911 = {1{`RANDOM}};
  px_buffer_455_g = _RAND_911[7:0];
  _RAND_912 = {1{`RANDOM}};
  px_buffer_456_r = _RAND_912[7:0];
  _RAND_913 = {1{`RANDOM}};
  px_buffer_456_g = _RAND_913[7:0];
  _RAND_914 = {1{`RANDOM}};
  px_buffer_457_r = _RAND_914[7:0];
  _RAND_915 = {1{`RANDOM}};
  px_buffer_457_g = _RAND_915[7:0];
  _RAND_916 = {1{`RANDOM}};
  px_buffer_458_r = _RAND_916[7:0];
  _RAND_917 = {1{`RANDOM}};
  px_buffer_458_g = _RAND_917[7:0];
  _RAND_918 = {1{`RANDOM}};
  px_buffer_459_r = _RAND_918[7:0];
  _RAND_919 = {1{`RANDOM}};
  px_buffer_459_g = _RAND_919[7:0];
  _RAND_920 = {1{`RANDOM}};
  px_buffer_460_r = _RAND_920[7:0];
  _RAND_921 = {1{`RANDOM}};
  px_buffer_460_g = _RAND_921[7:0];
  _RAND_922 = {1{`RANDOM}};
  px_buffer_461_r = _RAND_922[7:0];
  _RAND_923 = {1{`RANDOM}};
  px_buffer_461_g = _RAND_923[7:0];
  _RAND_924 = {1{`RANDOM}};
  px_buffer_462_r = _RAND_924[7:0];
  _RAND_925 = {1{`RANDOM}};
  px_buffer_462_g = _RAND_925[7:0];
  _RAND_926 = {1{`RANDOM}};
  px_buffer_463_r = _RAND_926[7:0];
  _RAND_927 = {1{`RANDOM}};
  px_buffer_463_g = _RAND_927[7:0];
  _RAND_928 = {1{`RANDOM}};
  px_buffer_464_r = _RAND_928[7:0];
  _RAND_929 = {1{`RANDOM}};
  px_buffer_464_g = _RAND_929[7:0];
  _RAND_930 = {1{`RANDOM}};
  px_buffer_465_r = _RAND_930[7:0];
  _RAND_931 = {1{`RANDOM}};
  px_buffer_465_g = _RAND_931[7:0];
  _RAND_932 = {1{`RANDOM}};
  px_buffer_466_r = _RAND_932[7:0];
  _RAND_933 = {1{`RANDOM}};
  px_buffer_466_g = _RAND_933[7:0];
  _RAND_934 = {1{`RANDOM}};
  px_buffer_467_r = _RAND_934[7:0];
  _RAND_935 = {1{`RANDOM}};
  px_buffer_467_g = _RAND_935[7:0];
  _RAND_936 = {1{`RANDOM}};
  px_buffer_468_r = _RAND_936[7:0];
  _RAND_937 = {1{`RANDOM}};
  px_buffer_468_g = _RAND_937[7:0];
  _RAND_938 = {1{`RANDOM}};
  px_buffer_469_r = _RAND_938[7:0];
  _RAND_939 = {1{`RANDOM}};
  px_buffer_469_g = _RAND_939[7:0];
  _RAND_940 = {1{`RANDOM}};
  px_buffer_470_r = _RAND_940[7:0];
  _RAND_941 = {1{`RANDOM}};
  px_buffer_470_g = _RAND_941[7:0];
  _RAND_942 = {1{`RANDOM}};
  px_buffer_471_r = _RAND_942[7:0];
  _RAND_943 = {1{`RANDOM}};
  px_buffer_471_g = _RAND_943[7:0];
  _RAND_944 = {1{`RANDOM}};
  px_buffer_472_r = _RAND_944[7:0];
  _RAND_945 = {1{`RANDOM}};
  px_buffer_472_g = _RAND_945[7:0];
  _RAND_946 = {1{`RANDOM}};
  px_buffer_473_r = _RAND_946[7:0];
  _RAND_947 = {1{`RANDOM}};
  px_buffer_473_g = _RAND_947[7:0];
  _RAND_948 = {1{`RANDOM}};
  px_buffer_474_r = _RAND_948[7:0];
  _RAND_949 = {1{`RANDOM}};
  px_buffer_474_g = _RAND_949[7:0];
  _RAND_950 = {1{`RANDOM}};
  px_buffer_475_r = _RAND_950[7:0];
  _RAND_951 = {1{`RANDOM}};
  px_buffer_475_g = _RAND_951[7:0];
  _RAND_952 = {1{`RANDOM}};
  px_buffer_476_r = _RAND_952[7:0];
  _RAND_953 = {1{`RANDOM}};
  px_buffer_476_g = _RAND_953[7:0];
  _RAND_954 = {1{`RANDOM}};
  px_buffer_477_r = _RAND_954[7:0];
  _RAND_955 = {1{`RANDOM}};
  px_buffer_477_g = _RAND_955[7:0];
  _RAND_956 = {1{`RANDOM}};
  px_buffer_478_r = _RAND_956[7:0];
  _RAND_957 = {1{`RANDOM}};
  px_buffer_478_g = _RAND_957[7:0];
  _RAND_958 = {1{`RANDOM}};
  px_buffer_479_r = _RAND_958[7:0];
  _RAND_959 = {1{`RANDOM}};
  px_buffer_479_g = _RAND_959[7:0];
  _RAND_960 = {1{`RANDOM}};
  px_buffer_480_r = _RAND_960[7:0];
  _RAND_961 = {1{`RANDOM}};
  px_buffer_480_g = _RAND_961[7:0];
  _RAND_962 = {1{`RANDOM}};
  px_buffer_481_r = _RAND_962[7:0];
  _RAND_963 = {1{`RANDOM}};
  px_buffer_481_g = _RAND_963[7:0];
  _RAND_964 = {1{`RANDOM}};
  px_buffer_482_r = _RAND_964[7:0];
  _RAND_965 = {1{`RANDOM}};
  px_buffer_482_g = _RAND_965[7:0];
  _RAND_966 = {1{`RANDOM}};
  px_buffer_483_r = _RAND_966[7:0];
  _RAND_967 = {1{`RANDOM}};
  px_buffer_483_g = _RAND_967[7:0];
  _RAND_968 = {1{`RANDOM}};
  px_buffer_484_r = _RAND_968[7:0];
  _RAND_969 = {1{`RANDOM}};
  px_buffer_484_g = _RAND_969[7:0];
  _RAND_970 = {1{`RANDOM}};
  px_buffer_485_r = _RAND_970[7:0];
  _RAND_971 = {1{`RANDOM}};
  px_buffer_485_g = _RAND_971[7:0];
  _RAND_972 = {1{`RANDOM}};
  px_buffer_486_r = _RAND_972[7:0];
  _RAND_973 = {1{`RANDOM}};
  px_buffer_486_g = _RAND_973[7:0];
  _RAND_974 = {1{`RANDOM}};
  px_buffer_487_r = _RAND_974[7:0];
  _RAND_975 = {1{`RANDOM}};
  px_buffer_487_g = _RAND_975[7:0];
  _RAND_976 = {1{`RANDOM}};
  px_buffer_488_r = _RAND_976[7:0];
  _RAND_977 = {1{`RANDOM}};
  px_buffer_488_g = _RAND_977[7:0];
  _RAND_978 = {1{`RANDOM}};
  px_buffer_489_r = _RAND_978[7:0];
  _RAND_979 = {1{`RANDOM}};
  px_buffer_489_g = _RAND_979[7:0];
  _RAND_980 = {1{`RANDOM}};
  px_buffer_490_r = _RAND_980[7:0];
  _RAND_981 = {1{`RANDOM}};
  px_buffer_490_g = _RAND_981[7:0];
  _RAND_982 = {1{`RANDOM}};
  px_buffer_491_r = _RAND_982[7:0];
  _RAND_983 = {1{`RANDOM}};
  px_buffer_491_g = _RAND_983[7:0];
  _RAND_984 = {1{`RANDOM}};
  px_buffer_492_r = _RAND_984[7:0];
  _RAND_985 = {1{`RANDOM}};
  px_buffer_492_g = _RAND_985[7:0];
  _RAND_986 = {1{`RANDOM}};
  px_buffer_493_r = _RAND_986[7:0];
  _RAND_987 = {1{`RANDOM}};
  px_buffer_493_g = _RAND_987[7:0];
  _RAND_988 = {1{`RANDOM}};
  px_buffer_494_r = _RAND_988[7:0];
  _RAND_989 = {1{`RANDOM}};
  px_buffer_494_g = _RAND_989[7:0];
  _RAND_990 = {1{`RANDOM}};
  px_buffer_495_r = _RAND_990[7:0];
  _RAND_991 = {1{`RANDOM}};
  px_buffer_495_g = _RAND_991[7:0];
  _RAND_992 = {1{`RANDOM}};
  px_buffer_496_r = _RAND_992[7:0];
  _RAND_993 = {1{`RANDOM}};
  px_buffer_496_g = _RAND_993[7:0];
  _RAND_994 = {1{`RANDOM}};
  px_buffer_497_r = _RAND_994[7:0];
  _RAND_995 = {1{`RANDOM}};
  px_buffer_497_g = _RAND_995[7:0];
  _RAND_996 = {1{`RANDOM}};
  px_buffer_498_r = _RAND_996[7:0];
  _RAND_997 = {1{`RANDOM}};
  px_buffer_498_g = _RAND_997[7:0];
  _RAND_998 = {1{`RANDOM}};
  px_buffer_499_r = _RAND_998[7:0];
  _RAND_999 = {1{`RANDOM}};
  px_buffer_499_g = _RAND_999[7:0];
  _RAND_1000 = {1{`RANDOM}};
  px_buffer_500_r = _RAND_1000[7:0];
  _RAND_1001 = {1{`RANDOM}};
  px_buffer_500_g = _RAND_1001[7:0];
  _RAND_1002 = {1{`RANDOM}};
  px_buffer_501_r = _RAND_1002[7:0];
  _RAND_1003 = {1{`RANDOM}};
  px_buffer_501_g = _RAND_1003[7:0];
  _RAND_1004 = {1{`RANDOM}};
  px_buffer_502_r = _RAND_1004[7:0];
  _RAND_1005 = {1{`RANDOM}};
  px_buffer_502_g = _RAND_1005[7:0];
  _RAND_1006 = {1{`RANDOM}};
  px_buffer_503_r = _RAND_1006[7:0];
  _RAND_1007 = {1{`RANDOM}};
  px_buffer_503_g = _RAND_1007[7:0];
  _RAND_1008 = {1{`RANDOM}};
  px_buffer_504_r = _RAND_1008[7:0];
  _RAND_1009 = {1{`RANDOM}};
  px_buffer_504_g = _RAND_1009[7:0];
  _RAND_1010 = {1{`RANDOM}};
  px_buffer_505_r = _RAND_1010[7:0];
  _RAND_1011 = {1{`RANDOM}};
  px_buffer_505_g = _RAND_1011[7:0];
  _RAND_1012 = {1{`RANDOM}};
  px_buffer_506_r = _RAND_1012[7:0];
  _RAND_1013 = {1{`RANDOM}};
  px_buffer_506_g = _RAND_1013[7:0];
  _RAND_1014 = {1{`RANDOM}};
  px_buffer_507_r = _RAND_1014[7:0];
  _RAND_1015 = {1{`RANDOM}};
  px_buffer_507_g = _RAND_1015[7:0];
  _RAND_1016 = {1{`RANDOM}};
  px_buffer_508_r = _RAND_1016[7:0];
  _RAND_1017 = {1{`RANDOM}};
  px_buffer_508_g = _RAND_1017[7:0];
  _RAND_1018 = {1{`RANDOM}};
  px_buffer_509_r = _RAND_1018[7:0];
  _RAND_1019 = {1{`RANDOM}};
  px_buffer_509_g = _RAND_1019[7:0];
  _RAND_1020 = {1{`RANDOM}};
  px_buffer_510_r = _RAND_1020[7:0];
  _RAND_1021 = {1{`RANDOM}};
  px_buffer_510_g = _RAND_1021[7:0];
  _RAND_1022 = {1{`RANDOM}};
  px_buffer_511_r = _RAND_1022[7:0];
  _RAND_1023 = {1{`RANDOM}};
  px_buffer_511_g = _RAND_1023[7:0];
  _RAND_1024 = {1{`RANDOM}};
  px_buffer_512_r = _RAND_1024[7:0];
  _RAND_1025 = {1{`RANDOM}};
  px_buffer_512_g = _RAND_1025[7:0];
  _RAND_1026 = {1{`RANDOM}};
  px_buffer_513_r = _RAND_1026[7:0];
  _RAND_1027 = {1{`RANDOM}};
  px_buffer_513_g = _RAND_1027[7:0];
  _RAND_1028 = {1{`RANDOM}};
  px_buffer_514_r = _RAND_1028[7:0];
  _RAND_1029 = {1{`RANDOM}};
  px_buffer_514_g = _RAND_1029[7:0];
  _RAND_1030 = {1{`RANDOM}};
  px_buffer_515_r = _RAND_1030[7:0];
  _RAND_1031 = {1{`RANDOM}};
  px_buffer_515_g = _RAND_1031[7:0];
  _RAND_1032 = {1{`RANDOM}};
  px_buffer_516_r = _RAND_1032[7:0];
  _RAND_1033 = {1{`RANDOM}};
  px_buffer_516_g = _RAND_1033[7:0];
  _RAND_1034 = {1{`RANDOM}};
  px_buffer_517_r = _RAND_1034[7:0];
  _RAND_1035 = {1{`RANDOM}};
  px_buffer_517_g = _RAND_1035[7:0];
  _RAND_1036 = {1{`RANDOM}};
  px_buffer_518_r = _RAND_1036[7:0];
  _RAND_1037 = {1{`RANDOM}};
  px_buffer_518_g = _RAND_1037[7:0];
  _RAND_1038 = {1{`RANDOM}};
  px_buffer_519_r = _RAND_1038[7:0];
  _RAND_1039 = {1{`RANDOM}};
  px_buffer_519_g = _RAND_1039[7:0];
  _RAND_1040 = {1{`RANDOM}};
  px_buffer_520_r = _RAND_1040[7:0];
  _RAND_1041 = {1{`RANDOM}};
  px_buffer_520_g = _RAND_1041[7:0];
  _RAND_1042 = {1{`RANDOM}};
  px_buffer_521_r = _RAND_1042[7:0];
  _RAND_1043 = {1{`RANDOM}};
  px_buffer_521_g = _RAND_1043[7:0];
  _RAND_1044 = {1{`RANDOM}};
  px_buffer_522_r = _RAND_1044[7:0];
  _RAND_1045 = {1{`RANDOM}};
  px_buffer_522_g = _RAND_1045[7:0];
  _RAND_1046 = {1{`RANDOM}};
  px_buffer_523_r = _RAND_1046[7:0];
  _RAND_1047 = {1{`RANDOM}};
  px_buffer_523_g = _RAND_1047[7:0];
  _RAND_1048 = {1{`RANDOM}};
  px_buffer_524_r = _RAND_1048[7:0];
  _RAND_1049 = {1{`RANDOM}};
  px_buffer_524_g = _RAND_1049[7:0];
  _RAND_1050 = {1{`RANDOM}};
  px_buffer_525_r = _RAND_1050[7:0];
  _RAND_1051 = {1{`RANDOM}};
  px_buffer_525_g = _RAND_1051[7:0];
  _RAND_1052 = {1{`RANDOM}};
  px_buffer_526_r = _RAND_1052[7:0];
  _RAND_1053 = {1{`RANDOM}};
  px_buffer_526_g = _RAND_1053[7:0];
  _RAND_1054 = {1{`RANDOM}};
  px_buffer_527_r = _RAND_1054[7:0];
  _RAND_1055 = {1{`RANDOM}};
  px_buffer_527_g = _RAND_1055[7:0];
  _RAND_1056 = {1{`RANDOM}};
  px_buffer_528_r = _RAND_1056[7:0];
  _RAND_1057 = {1{`RANDOM}};
  px_buffer_528_g = _RAND_1057[7:0];
  _RAND_1058 = {1{`RANDOM}};
  px_buffer_529_r = _RAND_1058[7:0];
  _RAND_1059 = {1{`RANDOM}};
  px_buffer_529_g = _RAND_1059[7:0];
  _RAND_1060 = {1{`RANDOM}};
  px_buffer_530_r = _RAND_1060[7:0];
  _RAND_1061 = {1{`RANDOM}};
  px_buffer_530_g = _RAND_1061[7:0];
  _RAND_1062 = {1{`RANDOM}};
  px_buffer_531_r = _RAND_1062[7:0];
  _RAND_1063 = {1{`RANDOM}};
  px_buffer_531_g = _RAND_1063[7:0];
  _RAND_1064 = {1{`RANDOM}};
  px_buffer_532_r = _RAND_1064[7:0];
  _RAND_1065 = {1{`RANDOM}};
  px_buffer_532_g = _RAND_1065[7:0];
  _RAND_1066 = {1{`RANDOM}};
  px_buffer_533_r = _RAND_1066[7:0];
  _RAND_1067 = {1{`RANDOM}};
  px_buffer_533_g = _RAND_1067[7:0];
  _RAND_1068 = {1{`RANDOM}};
  px_buffer_534_r = _RAND_1068[7:0];
  _RAND_1069 = {1{`RANDOM}};
  px_buffer_534_g = _RAND_1069[7:0];
  _RAND_1070 = {1{`RANDOM}};
  px_buffer_535_r = _RAND_1070[7:0];
  _RAND_1071 = {1{`RANDOM}};
  px_buffer_535_g = _RAND_1071[7:0];
  _RAND_1072 = {1{`RANDOM}};
  px_buffer_536_r = _RAND_1072[7:0];
  _RAND_1073 = {1{`RANDOM}};
  px_buffer_536_g = _RAND_1073[7:0];
  _RAND_1074 = {1{`RANDOM}};
  px_buffer_537_r = _RAND_1074[7:0];
  _RAND_1075 = {1{`RANDOM}};
  px_buffer_537_g = _RAND_1075[7:0];
  _RAND_1076 = {1{`RANDOM}};
  px_buffer_538_r = _RAND_1076[7:0];
  _RAND_1077 = {1{`RANDOM}};
  px_buffer_538_g = _RAND_1077[7:0];
  _RAND_1078 = {1{`RANDOM}};
  px_buffer_539_r = _RAND_1078[7:0];
  _RAND_1079 = {1{`RANDOM}};
  px_buffer_539_g = _RAND_1079[7:0];
  _RAND_1080 = {1{`RANDOM}};
  px_buffer_540_r = _RAND_1080[7:0];
  _RAND_1081 = {1{`RANDOM}};
  px_buffer_540_g = _RAND_1081[7:0];
  _RAND_1082 = {1{`RANDOM}};
  px_buffer_541_r = _RAND_1082[7:0];
  _RAND_1083 = {1{`RANDOM}};
  px_buffer_541_g = _RAND_1083[7:0];
  _RAND_1084 = {1{`RANDOM}};
  px_buffer_542_r = _RAND_1084[7:0];
  _RAND_1085 = {1{`RANDOM}};
  px_buffer_542_g = _RAND_1085[7:0];
  _RAND_1086 = {1{`RANDOM}};
  px_buffer_543_r = _RAND_1086[7:0];
  _RAND_1087 = {1{`RANDOM}};
  px_buffer_543_g = _RAND_1087[7:0];
  _RAND_1088 = {1{`RANDOM}};
  px_buffer_544_r = _RAND_1088[7:0];
  _RAND_1089 = {1{`RANDOM}};
  px_buffer_544_g = _RAND_1089[7:0];
  _RAND_1090 = {1{`RANDOM}};
  px_buffer_545_r = _RAND_1090[7:0];
  _RAND_1091 = {1{`RANDOM}};
  px_buffer_545_g = _RAND_1091[7:0];
  _RAND_1092 = {1{`RANDOM}};
  px_buffer_546_r = _RAND_1092[7:0];
  _RAND_1093 = {1{`RANDOM}};
  px_buffer_546_g = _RAND_1093[7:0];
  _RAND_1094 = {1{`RANDOM}};
  px_buffer_547_r = _RAND_1094[7:0];
  _RAND_1095 = {1{`RANDOM}};
  px_buffer_547_g = _RAND_1095[7:0];
  _RAND_1096 = {1{`RANDOM}};
  px_buffer_548_r = _RAND_1096[7:0];
  _RAND_1097 = {1{`RANDOM}};
  px_buffer_548_g = _RAND_1097[7:0];
  _RAND_1098 = {1{`RANDOM}};
  px_buffer_549_r = _RAND_1098[7:0];
  _RAND_1099 = {1{`RANDOM}};
  px_buffer_549_g = _RAND_1099[7:0];
  _RAND_1100 = {1{`RANDOM}};
  px_buffer_550_r = _RAND_1100[7:0];
  _RAND_1101 = {1{`RANDOM}};
  px_buffer_550_g = _RAND_1101[7:0];
  _RAND_1102 = {1{`RANDOM}};
  px_buffer_551_r = _RAND_1102[7:0];
  _RAND_1103 = {1{`RANDOM}};
  px_buffer_551_g = _RAND_1103[7:0];
  _RAND_1104 = {1{`RANDOM}};
  px_buffer_552_r = _RAND_1104[7:0];
  _RAND_1105 = {1{`RANDOM}};
  px_buffer_552_g = _RAND_1105[7:0];
  _RAND_1106 = {1{`RANDOM}};
  px_buffer_553_r = _RAND_1106[7:0];
  _RAND_1107 = {1{`RANDOM}};
  px_buffer_553_g = _RAND_1107[7:0];
  _RAND_1108 = {1{`RANDOM}};
  px_buffer_554_r = _RAND_1108[7:0];
  _RAND_1109 = {1{`RANDOM}};
  px_buffer_554_g = _RAND_1109[7:0];
  _RAND_1110 = {1{`RANDOM}};
  px_buffer_555_r = _RAND_1110[7:0];
  _RAND_1111 = {1{`RANDOM}};
  px_buffer_555_g = _RAND_1111[7:0];
  _RAND_1112 = {1{`RANDOM}};
  px_buffer_556_r = _RAND_1112[7:0];
  _RAND_1113 = {1{`RANDOM}};
  px_buffer_556_g = _RAND_1113[7:0];
  _RAND_1114 = {1{`RANDOM}};
  px_buffer_557_r = _RAND_1114[7:0];
  _RAND_1115 = {1{`RANDOM}};
  px_buffer_557_g = _RAND_1115[7:0];
  _RAND_1116 = {1{`RANDOM}};
  px_buffer_558_r = _RAND_1116[7:0];
  _RAND_1117 = {1{`RANDOM}};
  px_buffer_558_g = _RAND_1117[7:0];
  _RAND_1118 = {1{`RANDOM}};
  px_buffer_559_r = _RAND_1118[7:0];
  _RAND_1119 = {1{`RANDOM}};
  px_buffer_559_g = _RAND_1119[7:0];
  _RAND_1120 = {1{`RANDOM}};
  px_buffer_560_r = _RAND_1120[7:0];
  _RAND_1121 = {1{`RANDOM}};
  px_buffer_560_g = _RAND_1121[7:0];
  _RAND_1122 = {1{`RANDOM}};
  px_buffer_561_r = _RAND_1122[7:0];
  _RAND_1123 = {1{`RANDOM}};
  px_buffer_561_g = _RAND_1123[7:0];
  _RAND_1124 = {1{`RANDOM}};
  px_buffer_562_r = _RAND_1124[7:0];
  _RAND_1125 = {1{`RANDOM}};
  px_buffer_562_g = _RAND_1125[7:0];
  _RAND_1126 = {1{`RANDOM}};
  px_buffer_563_r = _RAND_1126[7:0];
  _RAND_1127 = {1{`RANDOM}};
  px_buffer_563_g = _RAND_1127[7:0];
  _RAND_1128 = {1{`RANDOM}};
  px_buffer_564_r = _RAND_1128[7:0];
  _RAND_1129 = {1{`RANDOM}};
  px_buffer_564_g = _RAND_1129[7:0];
  _RAND_1130 = {1{`RANDOM}};
  px_buffer_565_r = _RAND_1130[7:0];
  _RAND_1131 = {1{`RANDOM}};
  px_buffer_565_g = _RAND_1131[7:0];
  _RAND_1132 = {1{`RANDOM}};
  px_buffer_566_r = _RAND_1132[7:0];
  _RAND_1133 = {1{`RANDOM}};
  px_buffer_566_g = _RAND_1133[7:0];
  _RAND_1134 = {1{`RANDOM}};
  px_buffer_567_r = _RAND_1134[7:0];
  _RAND_1135 = {1{`RANDOM}};
  px_buffer_567_g = _RAND_1135[7:0];
  _RAND_1136 = {1{`RANDOM}};
  px_buffer_568_r = _RAND_1136[7:0];
  _RAND_1137 = {1{`RANDOM}};
  px_buffer_568_g = _RAND_1137[7:0];
  _RAND_1138 = {1{`RANDOM}};
  px_buffer_569_r = _RAND_1138[7:0];
  _RAND_1139 = {1{`RANDOM}};
  px_buffer_569_g = _RAND_1139[7:0];
  _RAND_1140 = {1{`RANDOM}};
  px_buffer_570_r = _RAND_1140[7:0];
  _RAND_1141 = {1{`RANDOM}};
  px_buffer_570_g = _RAND_1141[7:0];
  _RAND_1142 = {1{`RANDOM}};
  px_buffer_571_r = _RAND_1142[7:0];
  _RAND_1143 = {1{`RANDOM}};
  px_buffer_571_g = _RAND_1143[7:0];
  _RAND_1144 = {1{`RANDOM}};
  px_buffer_572_r = _RAND_1144[7:0];
  _RAND_1145 = {1{`RANDOM}};
  px_buffer_572_g = _RAND_1145[7:0];
  _RAND_1146 = {1{`RANDOM}};
  px_buffer_573_r = _RAND_1146[7:0];
  _RAND_1147 = {1{`RANDOM}};
  px_buffer_573_g = _RAND_1147[7:0];
  _RAND_1148 = {1{`RANDOM}};
  px_buffer_574_r = _RAND_1148[7:0];
  _RAND_1149 = {1{`RANDOM}};
  px_buffer_574_g = _RAND_1149[7:0];
  _RAND_1150 = {1{`RANDOM}};
  px_buffer_575_r = _RAND_1150[7:0];
  _RAND_1151 = {1{`RANDOM}};
  px_buffer_575_g = _RAND_1151[7:0];
  _RAND_1152 = {1{`RANDOM}};
  px_buffer_576_r = _RAND_1152[7:0];
  _RAND_1153 = {1{`RANDOM}};
  px_buffer_576_g = _RAND_1153[7:0];
  _RAND_1154 = {1{`RANDOM}};
  px_buffer_577_r = _RAND_1154[7:0];
  _RAND_1155 = {1{`RANDOM}};
  px_buffer_577_g = _RAND_1155[7:0];
  _RAND_1156 = {1{`RANDOM}};
  px_buffer_578_r = _RAND_1156[7:0];
  _RAND_1157 = {1{`RANDOM}};
  px_buffer_578_g = _RAND_1157[7:0];
  _RAND_1158 = {1{`RANDOM}};
  px_buffer_579_r = _RAND_1158[7:0];
  _RAND_1159 = {1{`RANDOM}};
  px_buffer_579_g = _RAND_1159[7:0];
  _RAND_1160 = {1{`RANDOM}};
  px_buffer_580_r = _RAND_1160[7:0];
  _RAND_1161 = {1{`RANDOM}};
  px_buffer_580_g = _RAND_1161[7:0];
  _RAND_1162 = {1{`RANDOM}};
  px_buffer_581_r = _RAND_1162[7:0];
  _RAND_1163 = {1{`RANDOM}};
  px_buffer_581_g = _RAND_1163[7:0];
  _RAND_1164 = {1{`RANDOM}};
  px_buffer_582_r = _RAND_1164[7:0];
  _RAND_1165 = {1{`RANDOM}};
  px_buffer_582_g = _RAND_1165[7:0];
  _RAND_1166 = {1{`RANDOM}};
  px_buffer_583_r = _RAND_1166[7:0];
  _RAND_1167 = {1{`RANDOM}};
  px_buffer_583_g = _RAND_1167[7:0];
  _RAND_1168 = {1{`RANDOM}};
  px_buffer_584_r = _RAND_1168[7:0];
  _RAND_1169 = {1{`RANDOM}};
  px_buffer_584_g = _RAND_1169[7:0];
  _RAND_1170 = {1{`RANDOM}};
  px_buffer_585_r = _RAND_1170[7:0];
  _RAND_1171 = {1{`RANDOM}};
  px_buffer_585_g = _RAND_1171[7:0];
  _RAND_1172 = {1{`RANDOM}};
  px_buffer_586_r = _RAND_1172[7:0];
  _RAND_1173 = {1{`RANDOM}};
  px_buffer_586_g = _RAND_1173[7:0];
  _RAND_1174 = {1{`RANDOM}};
  px_buffer_587_r = _RAND_1174[7:0];
  _RAND_1175 = {1{`RANDOM}};
  px_buffer_587_g = _RAND_1175[7:0];
  _RAND_1176 = {1{`RANDOM}};
  px_buffer_588_r = _RAND_1176[7:0];
  _RAND_1177 = {1{`RANDOM}};
  px_buffer_588_g = _RAND_1177[7:0];
  _RAND_1178 = {1{`RANDOM}};
  px_buffer_589_r = _RAND_1178[7:0];
  _RAND_1179 = {1{`RANDOM}};
  px_buffer_589_g = _RAND_1179[7:0];
  _RAND_1180 = {1{`RANDOM}};
  px_buffer_590_r = _RAND_1180[7:0];
  _RAND_1181 = {1{`RANDOM}};
  px_buffer_590_g = _RAND_1181[7:0];
  _RAND_1182 = {1{`RANDOM}};
  px_buffer_591_r = _RAND_1182[7:0];
  _RAND_1183 = {1{`RANDOM}};
  px_buffer_591_g = _RAND_1183[7:0];
  _RAND_1184 = {1{`RANDOM}};
  px_buffer_592_r = _RAND_1184[7:0];
  _RAND_1185 = {1{`RANDOM}};
  px_buffer_592_g = _RAND_1185[7:0];
  _RAND_1186 = {1{`RANDOM}};
  px_buffer_593_r = _RAND_1186[7:0];
  _RAND_1187 = {1{`RANDOM}};
  px_buffer_593_g = _RAND_1187[7:0];
  _RAND_1188 = {1{`RANDOM}};
  px_buffer_594_r = _RAND_1188[7:0];
  _RAND_1189 = {1{`RANDOM}};
  px_buffer_594_g = _RAND_1189[7:0];
  _RAND_1190 = {1{`RANDOM}};
  px_buffer_595_r = _RAND_1190[7:0];
  _RAND_1191 = {1{`RANDOM}};
  px_buffer_595_g = _RAND_1191[7:0];
  _RAND_1192 = {1{`RANDOM}};
  px_buffer_596_r = _RAND_1192[7:0];
  _RAND_1193 = {1{`RANDOM}};
  px_buffer_596_g = _RAND_1193[7:0];
  _RAND_1194 = {1{`RANDOM}};
  px_buffer_597_r = _RAND_1194[7:0];
  _RAND_1195 = {1{`RANDOM}};
  px_buffer_597_g = _RAND_1195[7:0];
  _RAND_1196 = {1{`RANDOM}};
  px_buffer_598_r = _RAND_1196[7:0];
  _RAND_1197 = {1{`RANDOM}};
  px_buffer_598_g = _RAND_1197[7:0];
  _RAND_1198 = {1{`RANDOM}};
  px_buffer_599_r = _RAND_1198[7:0];
  _RAND_1199 = {1{`RANDOM}};
  px_buffer_599_g = _RAND_1199[7:0];
  _RAND_1200 = {1{`RANDOM}};
  px_buffer_600_r = _RAND_1200[7:0];
  _RAND_1201 = {1{`RANDOM}};
  px_buffer_600_g = _RAND_1201[7:0];
  _RAND_1202 = {1{`RANDOM}};
  px_buffer_601_r = _RAND_1202[7:0];
  _RAND_1203 = {1{`RANDOM}};
  px_buffer_601_g = _RAND_1203[7:0];
  _RAND_1204 = {1{`RANDOM}};
  px_buffer_602_r = _RAND_1204[7:0];
  _RAND_1205 = {1{`RANDOM}};
  px_buffer_602_g = _RAND_1205[7:0];
  _RAND_1206 = {1{`RANDOM}};
  px_buffer_603_r = _RAND_1206[7:0];
  _RAND_1207 = {1{`RANDOM}};
  px_buffer_603_g = _RAND_1207[7:0];
  _RAND_1208 = {1{`RANDOM}};
  px_buffer_604_r = _RAND_1208[7:0];
  _RAND_1209 = {1{`RANDOM}};
  px_buffer_604_g = _RAND_1209[7:0];
  _RAND_1210 = {1{`RANDOM}};
  px_buffer_605_r = _RAND_1210[7:0];
  _RAND_1211 = {1{`RANDOM}};
  px_buffer_605_g = _RAND_1211[7:0];
  _RAND_1212 = {1{`RANDOM}};
  px_buffer_606_r = _RAND_1212[7:0];
  _RAND_1213 = {1{`RANDOM}};
  px_buffer_606_g = _RAND_1213[7:0];
  _RAND_1214 = {1{`RANDOM}};
  px_buffer_607_r = _RAND_1214[7:0];
  _RAND_1215 = {1{`RANDOM}};
  px_buffer_607_g = _RAND_1215[7:0];
  _RAND_1216 = {1{`RANDOM}};
  px_buffer_608_r = _RAND_1216[7:0];
  _RAND_1217 = {1{`RANDOM}};
  px_buffer_608_g = _RAND_1217[7:0];
  _RAND_1218 = {1{`RANDOM}};
  px_buffer_609_r = _RAND_1218[7:0];
  _RAND_1219 = {1{`RANDOM}};
  px_buffer_609_g = _RAND_1219[7:0];
  _RAND_1220 = {1{`RANDOM}};
  px_buffer_610_r = _RAND_1220[7:0];
  _RAND_1221 = {1{`RANDOM}};
  px_buffer_610_g = _RAND_1221[7:0];
  _RAND_1222 = {1{`RANDOM}};
  px_buffer_611_r = _RAND_1222[7:0];
  _RAND_1223 = {1{`RANDOM}};
  px_buffer_611_g = _RAND_1223[7:0];
  _RAND_1224 = {1{`RANDOM}};
  px_buffer_612_r = _RAND_1224[7:0];
  _RAND_1225 = {1{`RANDOM}};
  px_buffer_612_g = _RAND_1225[7:0];
  _RAND_1226 = {1{`RANDOM}};
  px_buffer_613_r = _RAND_1226[7:0];
  _RAND_1227 = {1{`RANDOM}};
  px_buffer_613_g = _RAND_1227[7:0];
  _RAND_1228 = {1{`RANDOM}};
  px_buffer_614_r = _RAND_1228[7:0];
  _RAND_1229 = {1{`RANDOM}};
  px_buffer_614_g = _RAND_1229[7:0];
  _RAND_1230 = {1{`RANDOM}};
  px_buffer_615_r = _RAND_1230[7:0];
  _RAND_1231 = {1{`RANDOM}};
  px_buffer_615_g = _RAND_1231[7:0];
  _RAND_1232 = {1{`RANDOM}};
  px_buffer_616_r = _RAND_1232[7:0];
  _RAND_1233 = {1{`RANDOM}};
  px_buffer_616_g = _RAND_1233[7:0];
  _RAND_1234 = {1{`RANDOM}};
  px_buffer_617_r = _RAND_1234[7:0];
  _RAND_1235 = {1{`RANDOM}};
  px_buffer_617_g = _RAND_1235[7:0];
  _RAND_1236 = {1{`RANDOM}};
  px_buffer_618_r = _RAND_1236[7:0];
  _RAND_1237 = {1{`RANDOM}};
  px_buffer_618_g = _RAND_1237[7:0];
  _RAND_1238 = {1{`RANDOM}};
  px_buffer_619_r = _RAND_1238[7:0];
  _RAND_1239 = {1{`RANDOM}};
  px_buffer_619_g = _RAND_1239[7:0];
  _RAND_1240 = {1{`RANDOM}};
  px_buffer_620_r = _RAND_1240[7:0];
  _RAND_1241 = {1{`RANDOM}};
  px_buffer_620_g = _RAND_1241[7:0];
  _RAND_1242 = {1{`RANDOM}};
  px_buffer_621_r = _RAND_1242[7:0];
  _RAND_1243 = {1{`RANDOM}};
  px_buffer_621_g = _RAND_1243[7:0];
  _RAND_1244 = {1{`RANDOM}};
  px_buffer_622_r = _RAND_1244[7:0];
  _RAND_1245 = {1{`RANDOM}};
  px_buffer_622_g = _RAND_1245[7:0];
  _RAND_1246 = {1{`RANDOM}};
  px_buffer_623_r = _RAND_1246[7:0];
  _RAND_1247 = {1{`RANDOM}};
  px_buffer_623_g = _RAND_1247[7:0];
  _RAND_1248 = {1{`RANDOM}};
  px_buffer_624_r = _RAND_1248[7:0];
  _RAND_1249 = {1{`RANDOM}};
  px_buffer_624_g = _RAND_1249[7:0];
  _RAND_1250 = {1{`RANDOM}};
  px_buffer_625_r = _RAND_1250[7:0];
  _RAND_1251 = {1{`RANDOM}};
  px_buffer_625_g = _RAND_1251[7:0];
  _RAND_1252 = {1{`RANDOM}};
  px_buffer_626_r = _RAND_1252[7:0];
  _RAND_1253 = {1{`RANDOM}};
  px_buffer_626_g = _RAND_1253[7:0];
  _RAND_1254 = {1{`RANDOM}};
  px_buffer_627_r = _RAND_1254[7:0];
  _RAND_1255 = {1{`RANDOM}};
  px_buffer_627_g = _RAND_1255[7:0];
  _RAND_1256 = {1{`RANDOM}};
  px_buffer_628_r = _RAND_1256[7:0];
  _RAND_1257 = {1{`RANDOM}};
  px_buffer_628_g = _RAND_1257[7:0];
  _RAND_1258 = {1{`RANDOM}};
  px_buffer_629_r = _RAND_1258[7:0];
  _RAND_1259 = {1{`RANDOM}};
  px_buffer_629_g = _RAND_1259[7:0];
  _RAND_1260 = {1{`RANDOM}};
  px_buffer_630_r = _RAND_1260[7:0];
  _RAND_1261 = {1{`RANDOM}};
  px_buffer_630_g = _RAND_1261[7:0];
  _RAND_1262 = {1{`RANDOM}};
  px_buffer_631_r = _RAND_1262[7:0];
  _RAND_1263 = {1{`RANDOM}};
  px_buffer_631_g = _RAND_1263[7:0];
  _RAND_1264 = {1{`RANDOM}};
  px_buffer_632_r = _RAND_1264[7:0];
  _RAND_1265 = {1{`RANDOM}};
  px_buffer_632_g = _RAND_1265[7:0];
  _RAND_1266 = {1{`RANDOM}};
  px_buffer_633_r = _RAND_1266[7:0];
  _RAND_1267 = {1{`RANDOM}};
  px_buffer_633_g = _RAND_1267[7:0];
  _RAND_1268 = {1{`RANDOM}};
  px_buffer_634_r = _RAND_1268[7:0];
  _RAND_1269 = {1{`RANDOM}};
  px_buffer_634_g = _RAND_1269[7:0];
  _RAND_1270 = {1{`RANDOM}};
  px_buffer_635_r = _RAND_1270[7:0];
  _RAND_1271 = {1{`RANDOM}};
  px_buffer_635_g = _RAND_1271[7:0];
  _RAND_1272 = {1{`RANDOM}};
  px_buffer_636_r = _RAND_1272[7:0];
  _RAND_1273 = {1{`RANDOM}};
  px_buffer_636_g = _RAND_1273[7:0];
  _RAND_1274 = {1{`RANDOM}};
  px_buffer_637_r = _RAND_1274[7:0];
  _RAND_1275 = {1{`RANDOM}};
  px_buffer_637_g = _RAND_1275[7:0];
  _RAND_1276 = {1{`RANDOM}};
  px_buffer_638_r = _RAND_1276[7:0];
  _RAND_1277 = {1{`RANDOM}};
  px_buffer_638_g = _RAND_1277[7:0];
  _RAND_1278 = {1{`RANDOM}};
  px_buffer_639_r = _RAND_1278[7:0];
  _RAND_1279 = {1{`RANDOM}};
  px_buffer_639_g = _RAND_1279[7:0];
  _RAND_1280 = {1{`RANDOM}};
  last_px_r = _RAND_1280[7:0];
  _RAND_1281 = {1{`RANDOM}};
  last_px_g = _RAND_1281[7:0];
  _RAND_1282 = {1{`RANDOM}};
  REG = _RAND_1282[8:0];
  _RAND_1283 = {1{`RANDOM}};
  REG_1 = _RAND_1283[8:0];
  _RAND_1284 = {1{`RANDOM}};
  REG_3 = _RAND_1284[8:0];
  _RAND_1285 = {1{`RANDOM}};
  REG_4 = _RAND_1285[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
