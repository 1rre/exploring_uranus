��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����յ����.7N�W]{�����<El���NҜ݋_t'_?x���9Fg��:_�Rd�H-ǏQ�w���+��оW0�C�+?Ǒ���{�Y�U��D��j>���Bc;�P%��^v��(��0�*S'W�&��[��qq�����'A�ꏤ��R���c~ố-0�C�O4� �`iY�g�2$��wA�
FI-71�W{���� C "A�e�OYS���M��� �p�������ƚ�p��C�>w���`_$�9�#��dOlB�"D+�Hvgws�s[���=)�y��S{tf;�A�Z�3!���>zu~�q,�!4��c��9!P���{D�����~:��XE��i�|����J��z�ў'���p��p&��[T�>9��0�s���+sA�:O�JE4K��S[������2V�Ed��z�]02�oi2��]�`�N���nt6���T�,g�T�s��(�'���s	7�W�u�"������@h��G��������ߤ_���S@W
�b��R"Y�^1zK~(��:����n�9�j5O6�O�R /�>]Nd0��C�'�9ȇ���$(���O0��V�<���*o�e@���L� &,��}���Υ��,�L�c2��_��A�v��g0[ۧ�^�#~Z<�wapH��P���SU'��#@���J�_��b�����
A��{D�b_�>���2C��Oq����i�2px�N�ގ��T���=��)d���
��� ��Q��]ŀs�8��B��CJo0U��0BRh�*P?���H�l��Sj�^]�Q��Oj�('�����|H@��]� ֫7���KV��'h�[lRl#y�i6	Rٿ�?y��Q����

K	=]�!�񀈬6����﫰Բ�W_bQ��\B3�i������L&�s��}'�)q�`��U�����W������ak��JR���i����hw	��	zB���CӸ�����o���\�Y�if-�J\`˂�zł����q�G�mu�cۂ�Hp��P�7�«�#2���rԅU�.I����.�&JZZ����H�j�Y�v�jO��`VS������T<��%H)�*l@�]����K��MP�������dg~/0��,ڴ��u�9����4b F�_���/e~O`�i��;�(}�8?N�Q�|� �:�d���
4�V��b_JIǻ �݈�NxT��ڵ��g���f�OH��J�ݸ*�����m"!��=N��3�ǒ�����E����;��Y�	]�Lꧧ����U��\d�B=r4+o�v��.o~�ޜje�
,�wv��)�ϭϭ�����V��q��m`s^Ƃj\_�ڢۯ��̭V�#��#U߹��9�ָ��6�{�� �ߣR�4��=F��u�~�u�key�
��*��:�L��=��'�_���?�A�e�R]�/$��UQXH�ڨ<mU�4��mh� k��m0�?���)`�>�r�	&��%�@�yM�����k�` ��+�+n�x����8����*���-px�yf�u��u~=�(�(#�	n�d.�ݣ͞����~:N$Ju���1��J5 �h�L�9������k�1�Gh(����/:�F���0H686�	h�����w���M�����\��JW�^n��B�+}�[{�a�R�x�OJ&w9�?nO�!�dI2[�b�!�S"�,Q���X|�����%]�RG�f}���W���)���S�ؙ
i�{�v%?X۟=?e;��I,}K�T[>^EI�ח<� *��A�I~
�M�J*q��ܰOAX���f����it=�bՠ�B&��e�! /M8�"v�P}� ��ֳ�|a(s��u[�+��9����|�@e�܉��o��;���s��1NJ�yY./�HyaG��Njt���R4�)\���s>[XK�9`@��I��퉖)+.���]���U�/��grqG��%�+�ף��z�tN99���%R'��h��ZF��[�������jV��<;�z��W+]g��G��ϩ�jl�+��SYz^�b��\	U_�I������� ݪ��cs�aPF����Q5��O��rnw���.���}�{��U����W>�����Ͼl���XĶ�ƺ9Sa�|��o��%n���%�E�.��^Xo2���Yϧ4>&|��)}gԱZz�b�W�z,�+��V�4�oVk��Dφ;�F%�����ߩ�TS&�busoN8����Lu�s�7��dq��k[U�R�c[JP�8�&9WTd���� ���X30��6���:!X�iu��Ҩ��d6-Mq�-ߎ}m���0�Z�HY)Ť.��ڇ�t<g�;�8A�j���;1�����䈧	�<>��ΨR��h�/��/��|�^��_�[�|qe`t
�~������`��P�q�9��������Ϛ�y��o�w� �}�B��t�#�"��*�c� �T)i鮂Z?ѕ�}U<��X�҈v���V�$�`��S�vw�]�䀨�+�	��U�o����G0x���y�{���; 2�Q�u��,|��?d�(ȹ֮��q���Ubi!&�r�� &�:q,���NA���	�?��,�Z _�X��g�9��?����4�lC_m��As�D��`�4�����\ѡ�2�wJ���u1��\#bV�o��aA���(��@�zE}��=����V�l�U�EL�8�K _�� '�CӶ���a��k	X�Ta�O�S�d�p�(��wpq (�N?Qr;����h����M��Gc3ѐV����	��jE�Eo�F	�����2�Ĺ���ߗ��CL�e�x<���S���:7R-�i���1�8��*���l�*�Ckrn^��z���+�����v��5��EqҮ�(L�|R0ݑh<ob�D���PF�Js�d3K�o~�c{ �g��L*�;~u��v�5���f��K�x��Cˁ����� .����+r����=k
�!_ �-����d���,��7�&���K�E�罃�Mg�81��CXT����N���� 7T�1��[�I��As�	C����SZ�H���� ��1�t2��>��B�����C��j�"2>�jmF(�i��g��(�9�>m)�1�żAF]׃�[�����g��u��^ �L�湘�V[*�%�JX����}�!V+S_@{
��	<$�� ���!@��2��j�1���-Ȱ��0Ǉ�t.���ŵ ��9���1��D�:�tWۧ;몵ٮ�}�6J�Ǵ�$�F�t����N��8���>��}7�Zc�Zl�W2���Nk_��a�D�q i���NY�6}w�<�vt`gŘ������_����*哎��Gl���������q��_`��
�G��G���`V������g�
��*����f)r\���؂)}���?,��Ў��b��W ���Q�|�R�S37e:|�W���Z��..H(G���ՆT˶1��9�� 2{T6nރ Ћ	gjQ,�{�J�9g����+5�!0s^�`#� �P��}~|a�Vw\�V�
����L�vfS�!|d��an����*�w�_PH�� q�5<i����UA�YG��v^�R�8�afZ�A }�~NB�ۏ�0@t���g_2ߌ����	�z`��	�+��i0�~�c�z��S1�بE����i�n�����b)g]�$I�}�3r>�z�mز�پ�m��KĲΫȝt��� JVy�慃nV��Dl��ۮ�ID�F��]6�[yH;���M�G{�UU�z�u�h,/�dp+�eЊ����UD���.G��٤��"q2��n�Z;Y�q��t>v����dS�M���9�1��b��B�?!ۂ~)ihO��ω�����x��O
i୿Sh�d���#P�H��R}��:9�u8h�Tf��;�g�"yR_'�w�wԘ��Z���݆��	j��tVHfv�q9�U�%��qLq!�Z���<-/,�?���x��}���&���+ Q���s���Y׈,!]��7���桿���9n�el�1�΃Lar	KE���Y��.$��EI&ݢZ�(�U�e����_s�J}�cʿ� ʽ�l*�|7r�{�>�.����%W���9�\�ݺ�g
�NE����.�]��"s-O�׆�����GH[�*��%{��TE��?�D�h��!ʬs����FK�����;|�#&uU�h6�Ȑ��Jq,��d~�Q|�W Uޖ��}(Wד�����|	���2G�;���e���V�dR��@��@\��*o^�+X�`H[,�>Ϣ��I*"����õ�Eؠ�$┼�-"�%Pj�*� P���ɋ?�pM+�����MW}h󾱕��� �
�|P<WrW��
}��,�t�>��!���a-e�a�i�zϱ���?L��6��a?�w�%�mO���&�u���Y4[fs.W��@/���&-�L'�U*��$4M�vf}UA1-)R�YY[��qĹ���|_���|2�w8E��Vc0�����k�\j�o�≖�SQ�6�P�ɾ���{�]�m
�=wIrc&�x]Ћs�bz:������P�>i������ ����k'�6-ɥ\�z.�� J��3Ԯ�nN���XԬ�|ɻ�*���#� ��;���t��"ffW��3��.C�S�?f����%8S�8\� V��@�[��cĻ��ҳ���
�2�C���yeo4(��|���䭚�l����D��@���]˛o'L����@��ԏ٨V|e;�@��m��-Z�ݶj�V\y���c�T���RTbǬ�[��ёE�/�X��i��.w�R���Ԧ�9d�ͻ�Um<-;1�J�/iW�+s�A9���V�y\��/�_fh�c<cW�m�����x8J���p����~�����_���a��÷���r�Ԭ�ywB��&�n�>e�y O�y�Zs���͖j�����⢧�!ZT�c��:~�ݳT�Wp�	\��i����n��Ł�����!'x̞�[���0�j)gH&M5��6�Ĉ ��i*7p�����~���%|ݲ����SWr�����0�C�A�ͦB�n7��cɡg\�āVb'*�F���c�D���*ڐ�eߑˇ,9�G-�U�@<�[���K54W�5l���1�B�;Z�zn?%�K�l4�&Ȥ�`�O���4�I5<�L��=��N�d?B����zͩ��z��$v"��*���K���"jƝ�d���,��C/��S�(|�;Ɠ�w[,��7C��ya�H��d���p�8���� ��0��A�B�P�񗊻��#+_��/y�(i����=�㒘
F�n�� ��⛋Oj�ߜ/��*`��T�3���S"b�a%���Ux}dBV�c	�>�j?�o�k�*[�7��'�`��VçΉ���}ٙ����g{�A���*5N�5k7�AJ�9�jf�E�J�n�m	��d'��Y���J���}g���i��2L��L��#���yp�x��J��W$�bJ��F%��x�h4�
)9�t$�j}�RiJ�[&�Xm���xo��Zmu��> 
`7���!cJ#g$�_�s`W
m��[s�/��V�"F+����SݥV�dM��p6ɶ���0�M!y��Ga�{��i�\!S0�i��L��+ĳ�x�4j�y#��x��+�X0��~pyon��5W	�t"�U1�D��؎�[l̎���b���˻^�uz�HI7��P:�W�30r�"�WAJg�N${s���<�8�{z]i�s�}��ݔ+�����؂g�'���Ը���/��N�;*��])M����sa8/sd�?z`��[=%iF2h�~Z�=N���8��\6��F#h1��V%s������u~�a7�o]Ɯ�l+�-&�n�s�Z���9̯���S�_�I�5�-�S��2l��p�G���Ӧ-k9U�hg�d��c,�����r"a��)�@�Z�DLK~ָ�b�p���#.3�1��8�w/_�|�B	UK����u�kF��+��\~t�p����t�_s9���z�y_��oU�K���`jƘG?m6>�.��S�[w���-�^)&�Z�6(|a��p��c8,
�e}~�b���~Mh R"��öm]#��=�vLh>t�ᑈ�z�9�ce�)t���oN1��|eY�C�[ �(�<X��,�%=G��Yi��>Q�ǖ�a
=��=�&Q�)|=�'!n�Y�5p�$�\
�N������_(��#����A��_��WcU�Ͷ\�~苾*�Kf���5�%�D����3���R:`�Ct�(�]K�R��)�;.%5�SMl�v��!
� �Lb���og`���b;j�FÏ4�a��0�_��2ʵ��TLOs�u��I 0���~�����Q,P���>X�g��[�KQG�Ѩ�\�;��x?5����Jw��5��9U�n��)�١�^%�A���mh[~U���̀�WT��|H���<>��odʏ^N-�M�Qe-���cS�{UɞTZ�y��:�Cs�6�gB��W�m<_Hs�(��@���H����U���C,[��|�����3���{
$Y>�H���ie����I0��:� �&�� bB�G�@�	<�2m�4{q�O�d�Ă\AJ��SG!�)ܴ�/Q�� �"�&���:	�|�Ԟc�"@�K�$�0C��j����]߁s���MI��d]��:#���bAF�@�jx~��!0͠�c<���zP%��M��i���;���26
$)�F�$A�� +���B|v�p�	�����[t~��#��fO,�ȥ���l�<��!뤎_�Z��k��Ķ��}����3V���/]��!�������Y��(���[0u�ZvU=�����}"x��eaT�F9�W��(��t�rB��r�EQ��3G�K�ve��n,R�8���#�cm��}
`�fh-��i$ͼ��P
r�87ut�����gٍ�����^�3����G��t�3iK�����X��zTڹ둌�C��k��2⓷���/҇}�E��#Z��w�^�yWV�9��{K�be}�0?�)����s��)���o��� �~#�����~J�B0����<85D8>!�6s&�F�\ߵ֢�l����t���T�f�r7�2Y���R0��G{�u�3����z��E�H	��Df�<�x��(���8��:2a�����t���h�QGm�Ի�K�F�j�O���QKu���/�H<J#PC<� �F��~�:< e��N�}�7��y���L�E�I�:�g2a`����M����pd�'�'�·�LE�ӧ�B�D�0WĢﺧp�\Z���E���Y�<`a���H��fdӡ�/��㮈����������wf��s�^df0�Ia�3Kk_r�(�)��(�4T��a��e�.ţ�Z��TO�m�0��ƈ���=dC��&��s�6�0+=�@��=���8� т\�=���d??�z妅�G�8[�O:���K^.�dV��v��8a��i�}�t�O�O?v7Y_�V}�u4d�璕ś�Ő�[d�v%V��Xש&�����S&�ɔ�Y�i���"�u\�%���k]� ���`gE����8��T�t�?@���>�h�j�W�B�j�kw��/RJ�FX�NvǊ�UM&��-p��8Œ�K��/X �i[���G�$1�f�� 7��8��E�~��B�
9�����Y��?lm�5����޽�gN�|0�6~�<��Q3�������)�A�_ę,�?��,����}'�Ibx�+M��$�����%�bFm���-�[��������5�z` �lK��hظל����jX|-YJ`�T�ǃq�#�vw�7�ӡ���Z��PK�������{6�w�z��%��k蠺���k ��T�TY���
	�ʒn�����l$�+���T����Q���`>�{KCr7�����z2ތ�ǻ�c�dW���g��,`��M6��78�rث�����4��<��oQ�1;߷���X���uND���4�!�*�g���lv/�BV]N��@b;��a���a��p��k?q�-,� �w�wak�`�
�`��d�0���?\�~\�(�-ۣ��,�U�v��Yae�u��*��F���@���W�|��#�xe�T�D�V�)Q���^!�G�;��&*ط�}�H�V�����X�aI�
h���� ���Si'+X"�.�$��bn^|w������V$;r0&�҈߆�	�����������׺{=0:h����L�
=h�@��Hs��3lP_��Z������{���3��ȴ�����r�R�Q;�pȽ��f�/�g�g?�^���N�W�[�E��&D=<"4�D]����� H*��O|�6r�G��;5���S�n�c������`�N��\֨5=�_���[Ă�Q�s�0q��f��e��< �|Ǽw(��Q�^�g��H��e�}����2����k�X�G/�pZ���e�l*�v^��ձU?نe�o�E�r����?`Q���jP��Jbvb�6.�@+*��)�ʼ�յ�5����2�=f�
K�˺0"\��.*�=P����)�7	��2����r��^v�4��a�F`.�i����{6[ֲ\������j�]�߀軪�����PJ��7lIC��Ŋ�2VH����$��+�ԸT�M ;F腧�<'�4�a�^&!�t�6�:T�X�ꏮ���+;��Q��
�3�G�s9�fh!�[��}��5)Nh.�$ލ���Ѱ������7�ᇁy�7���^<�FFX���X=zX7%��Kz+(���k3�E��f�1�o��c�AL�A[٪���7xJ�����|�\�f��`o0���̐��cNC'U�)��[�祕�7�|
�y�������= dzbX�ǐ�t�|Ѳ�G��8�C-0�w(e�~�0^
o�ntKYH�jx#�ҨG�.,��J��.l���|ee
hB�$�d���h*�+����������;�Qk'5+0XІ�+��lB�(�rF/��m$GyL2����-x7��� �������-p�=q� ��|��C�.v�{�O�Z��Ϯ���矛�>b+�X�����װ8�_q�1�!���g�a������-�7�m2lN3!��3{�c�B�dV��~G]��:�aG�7�u��Ύ����i������"W-~�SE���e$��+ʡ������W:��M�!��Z2٘��o�
�(�[&��dU�,���G?{W[>��i�U~T��:7!�}!;����6D[��M�qL4���;�A,�(%I�C�2A���i8B�Yqkk�c�.
O��pZ�ܨL���ޕ��=}�4蠑�ϨP�H�E�����i�R,��� ����L<h�;-}$B��1�f_G�6�q�ͥT�S�HR�Dk��"���v�U���Z�<��Rv��=31�h������1$w~�%����E���ˋ/�R�t/�(]�f��p*�a��;�&�{	�_J�L
�%4�9:66s����M����7���X֖�@�1a�ޙ�.~K*�����Щ?�o�{	��Pl�qxc1;�ǩ��_�փ7>l,�v,��}h��H����^N��!l��J��E�>s���%���;)�%j�C6�L�{#1;���}�sؑ���M76�tzu��
2FR~��s�$�m�����8�a$/x �8���P{��k�ɐ0B�1��Ò}L�(�{�{�&�޸��?+�.ľ����_����16�u�Cϑs��yS�N�w��dw[���N,�%��j�,�����F���d����?.|�AQ�5�½�E��^a��ܸ�wvܦ����5�3�+��V~�`O����8��G��
���
�Q�x#X9�S�we3�KL��T'�R���yp���>\��K,�w��"����(C��*�����̫y�宑�5����MK��̡J�IrP��Ngm�D+��by�1�_:Ea	W]�v~;�7�����(��G2BI�$�Z_M3�ey�Þ23��خ�G�vzj~���e�H��^�	juy��S?L�gYg6�Ȳ�-����{*����0��;��]���SJ8�9
�С�~�o�3j
JDwQ]���)(����pϐ������;�X�)~�F�� 2.5 ����Ӗ������f�X�٘��A�r��d�T�F��jRmG�8��k���$m�FE@S�C��(���gnln*�
��*�S3^/���۷���D����;�7C������|��6i��i�t�y0�f�_S�MQ�ȋ��0BF��OY�F4�H��N$5���U���4�g���� Š1�i$��e�V,���g��Z�YXщ���O�	� ��&�W���(�ˆ�l|t)���lg�Cn0��iJ�,�8;��S� �mh�ͯ�i傱7*9�����