��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��tsn@;��e� ��;~�X��$շ�,��m����p���M�P�L,Ld�Зؤ��1Ej�fz�v�ՐL�l�J�s�p�{t��Ҩ��k`���n(W��0D�%�`O�;��i�(��^���N?U����3�`�>���'x0��.|����������]��֌�6�-R��>��q	U�G��4K�b!p�����r����#pSl섋~�".Q�D�ر�G�| �5�I5`�Ycx����$b�C�������+����a'<5	�Rc���M2�.e$��KW9�;U�hb#�)gmc�	��]�~:��W�gV����Y�C5���=v��Pc�5���֟n��'FT�'�<E=Nl��1^;@��F�^����c�n?�m1/hW�����v	@���_�<�����p���n�:1*p�]5��-��Y"b��k��V����C\Z%�\��3)rtd~���>8����S�M��`�$�� ����Ĕ��s��\`ɪ�nD֜�2�%H��~���� �cx5�xJ�Vئ���e����T;W�9b.�]�����5e�<�upV���n�(�G���ɤ��F�� ``�O�+%�q&��yWsN�����X��6%C��ΪOơĕ��-Yb6%,־N7���:s�x}>��
��/�c��S
�s|E�7�R��|x�[�����M�3I؇�1s�[�dS�����\�<�*J+P@Y,C��I�C�������
r�G������,AI��#�
��5V&��<#E*}k������6�3$Y-���Ҋc��y�j�L�Z�7{�ٱ܄f�.��Z��Z��:���_�Q�_���`�?�����!�@���c�3&�M��3ު�1w��DD�'z**i�Sh�mdS��زa�5wV|�=�T@8�mѭ���cY��YΈ
�҃���I��C��Gf�Q�Un�}� �撌59�q�0�KŰ>Q�)��k�Yژ)s�=��l�5����5�\R�Au�V *�j6"���h�#�H��r���
}�0� �_��Z�sp�	Uʧ�������Z9e�$��3rKLy}����oUB{+3y��X�y�@���p�Ӧg��W<4;9�!��[�����J�R���`�A�Z���`���@���}��	�uRs-��~��~�@�����&X�6�FVڋ��X@�`L�`y���Y�;P���+���L"QM���m~�mC��y���(�;�Gqq�m����t�"X+5:޾A���o���Z��r:�^��7��	�%��\v��pԵ~�,�%�R8ؔEe��Գ'y��8�f��^�*���بN$oOX�'��|�g�̭@(�̄�*T}.V�a�ZȤ�wC
�z�~��|���=��J�m��bxBg NeN��q��*� <��'�n�>%�N��3���8�>����w!m�yD�AK}9@-'�F�$�7��X�Y_��%t�2-�)���q˻��5Y����@� �[I��n���.|l�����җ=i>ʕF:5;��w��I`�s�f��Ie��udK�����%�������;�F�{\Vھ���
G+rX�:�o�T�A��<Q%�b�Oǀ���>��Ϋ|r������}��ITe�b��F�c���A3����,_s9&�&�qH�f�A�,��fJ
��D�{��p�HYb�����) �xN}D{�mJ���;F�A'�ݪ��,�ohS(v�紃r|�����%�`�;y�Tq2./ؽbe���u=Ӵ���2�d�h�%��������c�eD�������W�jTZ��v &]ܤ�{������%���9X���� q��B�v9]���`_�IV�y�)t$g�!��d�\w:�.I�ћ�kɌ����<S���^H������$q�2hCe��:��Ԫp��E���H����}Y�������GO_D>���=8w�r>yި4wj�r4�o�ٌ7"��wT=y[h�	���X�����s`dX~��~Yh�:M�?����� 
�^�;�z9�s�*��'���!$3�~��*�U6^4v@D��Վ�� ?a�)*�F�u�1ӧ�H��L�![�b���*N�ZG+���mM0���jCz�C��~�k���عL%��(��x�m���7�8�B�?z�ěf�VRJؐ� �Z��=i�`q�ܐ��������gg�|#u���j����q���n�d�b:��:���Lر��`�'����A&���>��b�?	��8љ�H�\��W�?��&	�"���YG�y}هOu'#5��͌ew�'�p��&5R]�3���y|��d�ִ�m�&��=�3��2Eut�,�D��5��UCб�z}+b�snkE)�Y��9�9������L�K��[)_��#��)����|�>x�"�wF�C�C�$���� �ٲ4B�*�m�l��Ѷ/Q&���+��'��]mJ0a����� 8r^m�|*�'��E��?ۙ��]|�>/n��?Kdn��i\g�JT�[aE
4��H|8��R���]C���}���0���WԍJg/0v�;R�w�3j)�p��� J��+Ǿ�CZ�D9�2	�	^��UD�T�kH
y܄J�ͷ�!M�9��w�ܘK��hBn� PT����Kء+�=��C|�FIĹw=����=�b\��e�wks��sr�ƴ蔊+�!�o�4�dT=m��&Cj��K�:��%+������&�),TQ�5{w�>FX1cS�rt%^}�7P����^�¡�̿�Y�2�MP���yٷ�L���������,-7�B��Nm���.�^T$"�詰��sh�ne:�̿��[���k�� \W���`��ܗ%�)�K�� 4���<(s!�����h��AJ��Â5Z���Ĺf&Ʃu�4ͺ�eO-ɐSY�տ�jmO��d�]B �r~�g=���i���L�rf*oJnh��W��<��H��V�Vcz��}-\Qƽ�C����D|D�J,�d^��d��u8'`�#�'�_?�Gyj�l���أ6M�7�&:��x)��C/��f�?f4]�>pi��H|�z���e�t�+@9�us�ߙ
c�UF<H�E��>~�-Nst^d��"|Aj�����4!� �B?�6l&LMLk*A�g��B0&���PΥf4G���%�{`,���燥d�X�������_V1*�.�z�+:2�m�����v�%��1l�B��'���b:;�j���xV� ʵ��N�FW@>��'�ŇdXY���� �_km�娮�ccP ĞQxTܻ:���R����;�#|��]����7q�y�|ׯ����q{���iW�X����a������tX$�6QO���$	�(A�\�羠��֕��$���}'V�/�ikpB�n�K�;OQ��W�)����f���Kb2�,a�%�,1fcÉ%�LM����9N�
��>��(��CT?�M��00����;y�m�N��QU�z��c�VU�й<�ǒ�ϐ=]g���Ʀv���΄g��q	�gX(/N�I��8Z�@J��D=py�s��QI�ͣ�f�ȏ˰g�d�S
�Ny�=*��WZD�1���T������#��Ac��O�M ~���q���Y�~�-����-�G���Vߘ�mtp��dU`�.R���I����TXB8W��E4�ʨ�^p]�\��,1쒴`R����9e�����'�"v4�o��Z����H!CZ�'���
���5{Ӫ	-�i L�����6�X]�����G%!��*ɁL��.JB��y����
�uMG�����ļD�X*�����"[���9�r̽�V/x��m���(f���W�	͏&��o�JIFs�&�Q�xەx��Nϙ