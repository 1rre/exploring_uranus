��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!� 7lw�9��:�6I0n��(Z���\��;��ݟ�f3Q#�Cݹl�X�j��Kd�ŗϨ����a;H\�&����P�p�V���R+ň���&�n�򖞘��ŧ4��@�S1��Y4�fR�Uig"X�?��"���n$��|��Ǘ�;}�)x�I��M;;����<�2Ķ�L�9p���[��tKJU��H����s�ܥ/lB�۲.gU�A\�4U��k���헧�bT�,���N��RʞO�BD�Ɓ�ͧ�f�䓵c ��'#u��K=�E��hѥ�Ȉ�x9N>�B�M �q%������_�m�1�75��3�&QnFK�İ��/�]W*��Q�-,�ݳ#;֌����G��q�?x�\]�)������ #1�sF�9�M�Á�f��I!��TL��8�e7�w~���X��GRl�w�nH��mi�V�?�U�a�t[��@��F/I����%����u�~#���]y;�'��@�ڠۗ��R���l��'E+N_t��^�-|5�^���޴F�:<LA�v��K���Z�f�`yb\�Gh㦉����
 �`v[��c���ķ+O;F'�rT�F���ݬ���jo�-��>��Ƌb��W�.�ƌ�,���&�L;����BY�Z�.��Mݩ�>��G��d��u5��k�P�~xK{�r�Ǆ�-��Q���*u΍<)�CȘ�d}�Y�~���cB=����`Z�0
3v���ql-��^#�p�,���ʒ+�W�C�kf�2�-���*�Pi�+H<��\���F%�1���}A7�QZ�f�(�||))�$Su1�ʠ���[Y�)x5O�'��+��-}�b�;MVJ�gg��;������5\����Ie��Ҕ`3�0�s$F7�+�L����n��v,c�z���YW'Q\��W$�'�ċ�ıT%����V� ���<:ǐ'K�.���[C��3����d5�X��Z?� I����B���N��u�/ç�]����0r�zi7�q�8��R�A��� ���rǆ%��}e����U�=��U��v�1]/t]A�\W�D��P��:�E�$�v�j��e��c,S��d���[�ΎY'�s�}�fޡb)I:���2c����W¯]��ߗPx�bi���}i��(��?���ݡ���+���9���w�澌q�����e���S$�­�*&&{�7L���P�ّUW�e�/�΃�O9O�o���{���S��^��'@N^�ϙ��vC�H�5CPmDI��v�!f^��%�6!�[̎�'ne��J��0{��@Њ�ڋ�Q��=D,���p��:�P��"�l\��DL�MOQ�+��t������m}Q�-vC~D��6>�&m�a��9�mO�R��l.[���V+M�V{��1����a<l�F�|��� ��� p3�����W�hLV�,W��³:,�ba�Jy���#�-%E�8��b�a�x�*$������P��0���L��ͨ��(i_��:�a�(���\}/��%�(��0���$����,\���S_9�^5͚r��p�~��r8G[+Y��K$�W#�&s�ޛU����Nb�H%��Ç�ΛX�^���"���N^��_��O�f[����y�W�$�0�����='oc2Py!�^\.��ڄ��V.��"��!��5V/M��(��y�[t�E}��*Y�C泜�T;V*g9�g�B��A�C�V��/O�6�|ԫ Q����js�l�&���H;�U&�bC�m��D��Ŕ�h�Ŵ��E�QS�2-����g,�;&ۃ?p9��� j��~�>�/�Z&�R(|"U�`"w�ߓG�QѐBq�zJ?E3��UŽ�
�vj/,W��6ɯˏ�lM�^��P"�~��Z�m���4��>ԋ��(�0�8�oS�j��=&k��at��X
c�L���������>�B£�x�h�4u(�I}#�D�H�w�U?2�a�Q����{���+��z)�\��=M��X�g�v��U���rb����伺��n{w�;��(����Д��C�~��)A��:)��\��� �2�mmC\��M��]R���=�
��O��QI[U�o��22�m��F��9
���nȲ��Ȝ��&����%X��  ��.����p�`�[���/���93����Z1��*�u\� |��]᧖-���
̯�P#5�I�W��N��"h�E���i��;�)��D��k�k�KkV]1ؾ�$IV3,��}O�y�z��_A����>��I�k
q�!U�)B�/��,HXb�ik&��y��s�%�5/�;�ό=�L2�L��7I!�p/2>��D�ꞽ
LY��Q�jiK[9� ����4S޴��`�`��vt�qE_o�%���Mr��x0Y�:.D��,�U�W�A��Iي�vw>7H<wi�~wB���ݫ�r_�u�sE�c��,�8���>�f
�PV�`�J���;�|��wnyz�qc����h�<m��r�k#���y�sۍc���	9Ğ����2@T'3mo@�/�K�<����d �+�������5b
�i�B(~�/��N�`B\�5��wNэ���k��	.e$?��o3�-1�x���Z=�fY�e�9�'�	�P���"��:U�3�n1xǆ5�� 3h�|qg%e��m�F�	,m>�d�uϘJ=C�ho��5��\^2�č�/�y�Eqv~�K��~�� Ix�(�&ǆ���_y..qQ>�$��ѹ��VgD 4���/G���ѫvnF����?��͠���ko�M�@�3�����69=�'��"n��4ð���[Gч�š�4�ނ��ׇ_�n�ջ�ѷ�/�?���.-�+��<�Vϝ�(�pX��b*ٺ:�%���+��h4�(�_u�-W�4��P������0�����OVa��"*԰٫1�b�S�B��t�UGγ1E@#��\	*֜6�$gִ���&J�I?E(D�~�Sy��,��&4w�d4,��+��H]�e��HaTt�R���i���Dp�?� ���֊w\P�{���m2�P�,�3Fº±Q�{���|��X��A��+�1�&*�o6����[R��N����`�O��K����/�����l�.�U��,�}��|�E�C+Ǳ�Q����ͱ�j6��:�,Ղ�E�O`TM���F�ߧEA�ӻ����w�;��q�M)�lz��s�Sb��o%=�.l����V�%�3YZ	�	�i��t^�n&S�pG�xb��3��������;�ۗ� ��S��&m*�F:ߣHW9�OW�a=�E�����k-&���V}|
8~��儉�s<��yz
[B��%�-���,�f��40an`WK*k"���d=V�go/���fBP �M�{�*������LI'��I={�$�h���4ǂ�e���޺9��kn;����HL��L��s�ةW��s@L�;�����5��P�j�V���׽c>�z�
��"vyW�rh�ƣ���.Ԙ࿰���V�g�1���!�$1ا��R�q��|������o�T9b�7w����ɬ��C<�X޸�m����C��i���P��*U�b([2��uY��M@��r��?듚�6�������z��"I.���:봜�����J�����~�#�߫��L^ �D1G_�R����k�g��S����*�!�P�E;�.�4��koh�y�%��p�aj!�o�t�F\��z���h�7ٓ�Ug.�����E�~�����k�����@�2������$g�QҚ������_�'���c�FQ
_�߇�@Ub��dĲ�]O��b�z����s蔰7����d�8�Y����kݷM�M<b�z�l����*�[�I�˜P�^C��h;؄oZ�MI5r������1{ď��~�ԣ�6�3�k'A�KK��-!k�~��kWc���_q��q��?�<��|�1�;mɦ��iB��$�Nj�'��Ͷ�2E5��@.=6�R����t�x/���$G\O�N5��B��\���/�ƘQ+����m�f�+�n�q��*:>/�	��5ǳ�M�VTi���)O�����-~k&9�Y�f�`���)!$��m��?�ǘ�4\�3u���CK3;� �h���8��kl�d��["�����&���%d,����Nz��@GbLw BV�vk���7f��/��#�NC>�~�PND��2�
.ȋ�y �&��Ͼ��އr�U��r��A�ci�i��q�/4�I Gܜ�F�՛]�*�E�Ɣ4,!J�+T������*����ۣ�<��o��U�-�����$��Wm�0t'x��/���_��JفhUS1����g�_�g����t�wu��@7�v�oLb=���n_{ED���A�*r�e���Ƥ�2���$Z5��N��mOX0�#�@x��*#��D�jf��̱z�������F�e̲8\���]�U?ik�(�f�?�}j͘�%W�����Q�e5f�ERx�h��=|��p�*�M�.����3a ����E*��;�j3r��b��ߧ3d�K���R�Y����R����i��J��S��?{j��Cf:��Z�2���~"��D%����Bk!$#N_9k�NS �)�`�Fb,R� ɓ�����L3��I���q3(���zO;̦qt]�Q�{���" /v��	�cNC+�{j9����s�]���+o,�&��r�F��5ۄI� �e9��̱0}�:����fo����5_.h���]ok�U�C�q ���1���i����~x���/$�p��j�*�_�s�F�����uY��q	p@˺}z&p�k� ���� �.ϛ1��S�&�o��"���uO�&�:rL���ƀ-|�)��5S�#���ۗG5��k1���"e���T�Wl~��&n�}|G�>[�6.v���H-��7d�8o_*	���#�����hGq��-�oI8>�j�S�3��N��6��8��N���E�����F��!���s��; ��� ���,X���e�%]=��� v׷{	�8�9�p! $��7+�1Q�x�of}�M)GW�J���se�C�脰�;7;�$��a8ִF���'��/>O����}�X�)t5����!F�7ۋ�2��D�L��`C�B{̃~ª&ɖ���EY1�c�eL��P�
9�d��(D��n9�韏UTF������ �V ��
����m�6�NZ�4���W6�d4ն����5�C�,���#�FD}�Q63�K�S\~�37K�� ~rV2!S�*v쁃�˔6��|c��ن��ߏT̝��o��JR����.����{���Df���:3\�H�7H{�
*I��J����a������*ȗi�Ғ���2�f���vR�yM�X�΁�go)�Qw����`Hd���^�r1�*�n�}R��&'�~_謮ZJ7*}���gE���$d��C��Ņ�WC!��ʷ���g.�b��(�Vm�8w�h�p�VEt�K_��%:���itʗ��#p�����tVAz�xJ�j �i��L҇�фb��-��D�@*�{�X�J�m�ϑ�wJ�"��kN��isS�!X�@kn}�C��$Y#=ud�=v�@�P
�P�[��j)ۜ�3O�v �4�Cz2��iGg{\q�P�q�H���^�w�I����(}кC�;!m�`��EfN�7x�>��z����N�tZ4�sUB�NI�
ps��q�v�XdS����Y�!mj�_�_�����o�Ou�o�kG��|z�GlcN�2�B�Zݵ��k�+�T�@i��d����5�Fj���>��q���W);z��~hFi�	�>��ޭAB�l�)�(0����Z�������~aV���s�RH���{�aX�߹��.�:�.��#o�MA�]q�HX.�r��h��h�:��r���NBԹn�Y���5�q8�hO[\j�jȀR��<|�r p���@��6�B7k�V��y�f
�_���M��3 �	��ޛ��.��Y(�.�V�I�6�C.x���Ĺ��6�9b�'�sZoh�d���sW�y��S�v�:��s �J��i�<��L���U�_��T��)� 5����ܶ�!X~�Dӫy�~���J.�0��ɞ�AN5�W�8�X��9��{���������FF����K
@���!9Z";k�hJ>Z�1�����'ߝo�_6��nW��V\���ᮓ+dd��KE	8�jAu'�m63�cϹ�?�E�����T�jt7�	���G�e�ެ��$�#iM^���Q�)�"��ͬ����\-u.�d#��=�W��9x�Cߓ�Q匆�(qC1ߜ�|���P����eU����6qG�������e������E��82]<���#"���ְ�&ˬ��g+�H��-��[N$^�'s=�����1��bH�����O���$΂�:�r�g�U)l'>���I��k�4��, ����neK���	¼��\�j�m�m�	mr���|��~��^��8���O)C>8�w'ZL�Q+��TCfz�э���V��q�j��{�p�n�Q�K�p�s��TtNO����9�;.i܂�FT�n1�'G�{i�c��]�ﬓ��_�	⣿:��J�ug��j����l-�2z�O=�������g��{�R�L�Y�BwD� ���1�KB�xi�]��R��&�"���Gr�nh���E�*s��yK]�q�w��Hn��>����<�z�׸i7��QI�O\cSs���g����2^��*Q��pn3;��@h䫖���a�d+ �J��^,|�k+A{ғ��c^0�^z�2�׸��9���A}Q!"tV���E�삜;�J��ț�Il�
-�����o]���'��d/����~;��kaw�+b���������"c�]�g�p¼U��V��Ϡ��Ѧ�W�GzPM\�f�2���,����(�4����Fq���4�M-#�N��bo˘h��M�r]q��	\êVj~g!r�~e�������
��