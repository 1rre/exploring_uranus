��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;������_$g��h��������"$��t�a�w~_�#��J�� 6:<�#T)��MqJ���K��� �Mv�:) GBNak���$8H�;��Ť_��I�'X=5Iټ
��2&�mn#=�y$\�L^um`E��\8[��`���dg�ދ�������DN�$	�F/���\������&�J�T	0�EC�Zg>���?� ��K��T��@6j&��I�8�ǭ�7��YE'����2'��]/��IB1p��"���l����b��d�yImd<2�אm���[��'Ӧl/��Jָ}��yn��s���vˆ�;�"����Ī�_X)��,����
�֣c誢$���������i�^C�!<ƅ�E��鍸j
Fl���e"iq8���_�_c�;a��֕�wؿ���p�?��TdW���c�{j��RM0��(OTz*��Cg���:��mŎ�N{0�QK�����%���ٛ��wT��0e���e������c�&ZH�sLXy�h��2ķ�=���!�܇+Y��).���QD]�1�i������j�Q\�t=hī���rZ�e�Ȩ�L��$g��a��ޅ 4"U�߲�����9�����fl��6�^pA���O�Ȍӏ%d���QtP��ٓ��Z�d����t#큮@�4b���P�Q1�����v��X��c�3�Pǒ��p?����!�w�һj�?��J�P�T�����Sr��?	jZ�#PM���	���L�q��kǠ��>S��m��CI̴�}ѕ>��E�)�@�'�ε�#x���I;]D_"���UY���f
N�j�0��TO:�vnҎ\N9�fl�4Vp{�Ϻ��1�}���%u�f�{����>�	 *g��JI��:�B�lIT�j+v�	�F>�����<�!��/q���a�]ۤ�YA���u�-�A��%�Z���3�&ie��G�S_�v8�D��P!������yG�T�4%��X�x��;��|[�2
TSh#���Wl/�(Ɇ,ܠ�xN��&q�ϋ2��#\��������htiK�kk���>�+{�Mh�F�Cx���0�5m(	�(�n��
��Y���61v�>k�_E���߲$�Z�5w�-0I,���7�0o�ě�B�|��n��f��a	�n�B�/�*��>4�7���]4䩔���`c������ư�b\�7��m3���\~���>J�ks�g��I���-��vY�K{�#�-�t��UWiU�ҟ�et|���Y��Ǵ�m��.�Oi����3��uc�|9l)Ǎ'�>��?������j(D)F�PS���!BE���G�����`��_�����E��_5#0��t�*�2��!��l���}��n�N���h�\o���(�P�(8�����z��.X�^ژ��/={/��h�`�i�y����7�s�-8� fau��B�g�x�6�Q���ニtn��ݦ�}�lu�}��`�
x.�O�Lݲ�YujIr�0����""�*čH�~Ah�.]�>�y���k]S�fw��ވ�l-;�W ���S��/Y�Y3��� �S�����M˳�I�-q��UE�A�T���J"H�3R=�c��U�I��S��֟���4jV�,�i�q��I;1S{�Fی�5	��ʳԞ��㝄{�_>�w��,�*�`��-KJ�B�]��	yX���i�U���;is�y\r���� �48����ЈM�� ����,2�͹�jO��$p:��؈(���x��A��Z8+�,��}"�39�Ql�d��!È�+�G� �L��B���.�i�}""c'Oo!�(��i�쯱Z�H9B���c�Oԕ"�`S���Cw��uaQ�Y��hO.`���p�1����✅U^)�J	s���}��m�΍��q�u���RG]�
��!�ݫBm/��yz�4���Cߦ���~��4�ʮ�b�L��{,���gI�#Qa!�����9����ڍ/�p�~��׳��b0w�6�5�釈0tr��dP������z���7%�گ�����2a�����n�\XѴ��L"r�#�{a���B�1��WT��c�� �ey%��W�������״E���I/<u�[�n����:�Ɨ��q���d�ˇr�x���6z��a
�P������ZE|L�]�8��� �������������3l��.@{[�7_˨�'��?�����njD���]�ǖU�׾����V�3g�WVb�M��k�1�sW��'ϒ�U�t5i(ɧL,/��L�Ή@�畧�{d�S�G񕀊��R'˪G�.���X�oS�Ǵ^j��\�O��8vq�^�b�ad
�{�G".����
#)�S��m��������όI�\0�5�]_��v��>�&�9I��n��Q� �Oe�̝�\�������~\�̈L/����w�z^��Hmw<�s��xM����x����J�f��I��P�Ԙa7�(���Մ�u�W��r���sm��=0�ҭz;�6<�/"�����<ϕ�fBX�9�F���W6��5����4���f���v�j_�|�&�_��F�6όu��Xo�dAr�b �},~r�pt�FX�g:(4ȵם�KOH�� sP���}��6/��A�	G�Ls�� .��u�� F��y�ׁ���DbJ*
j�,h �U���ߒN�n;r�gHc��x�a�����qq`1}�q3�L�1��|Y�|-�Ѐ1�T �����΁�ꔇ�|�N�ܻ6�,۲xS�V3S����|�o�(Wf|bȘ�'q�3#���Hl#�H�'��-(������Uۀg�u WQV�9���qa�� N��`W����2�7��S=^{�% !�Ԛu*�p���1g�n`�*y7���wA���{ʘ�-[�k.�	�������׶qkfI�"�z��3�vCI�����Or,�4�>hk��R��Uq�P��(�"�g���Y#s�
�����嗄Q�����<?E����|O6�$s�#��^�:�4�yʃ�O�x��&r��}�̾��ura۝�6�sG~�)��B��4���nL.�
��7�nA��j�ZE/.���R�A��"innm�`����ڙ𰋽�Y�M ρx< ���{�=���m���i�>�e$�g�	!��l)@���+o]�H3���Qe�i���S�4�?z]-N���[�Z��,C:���N֍Y�Q��z<|�-���2�B˛����_����U�c|Vrf���8��?<��6��1Y���X�0'oQ�2v���I?��5ʉN����>�.-���E;����C6�xŀ��:��@�.�41r/���wL�o�r`�[��[���]:0������F.�Cam��),� s�D�m��:�֙d������o��:�`t�0%2�w_�L�.( �i��k�j4�g�|Qa���&�,7DN�,�9�̍�S*�v�M��x�2$�|�"_��BU����tJ���wx�-�{a�b�V��S��jw/�K�G���\��L��,a�\�p�K�F�l����q+�Fk`�q�a$�T�H�%D4[��+$�7뱢��
���9��y ��a9��ʿGq��5 t�	�D$�[���ǻk��(�)���,���r��@Q>��b��Ϻ��M���xی���Y���G��fJ��q�eM���o�;�)�F��-$��]�����wQdl�̥�!T�������˘�{��x�mY�����c$ȣQ꾘�\�u�390��~�~3�T�S/�6��~R�ܾ}�>��MUl��	�{�X��,��?�]�1} �b\�/��T����T���l=(��>��v!��n�G�r'�դ�z��2,;K��o�	���rC�bD�m�����b-��;srKg=�Цe	O��y��$8�O:~�����|���c�=:T�q�H��һ^q����8����Ř���UάS�V+�{������k�j���Ȋ��U�����K�ph����𸡸�[L`��U)�H���U�t**��S��T��~Q7�ʰ��%vj���_��_ ����[{��4n���/% y��#�_:�U�� �N�0�P�"ʺ$��(��mp
����KtpQ�v��?�^6�SqjƑ�oV|����5�kJk>/�O�=��T:%�����ؓO��'�ut��}����eҘf��rE��>~4�(wo�g�ȧ���&&�&��qlAw�ǭ�v�W+���� C���Mv�� ʢ�/П����}�R7D0׌�O[ri��i.���NNn�#g,�c��������SM���h	3���epoo\�3o'�AH_��J:��Lj�%��(&zŶ�;��$t������I1����I�X�������:W���`����RU:qp�nZ�;�ulbN��y�o�,�g����|v���ȅ��mZ�>cl�G�%�*�k0�������5���R��I��� 4�����o������$���&/��Y�t��n�s����:�Fm���b��<�C� �%��^�%޸��;~�J��:�;��T�Qu�[�����ߕ�a�"+ �O�-�l��Z�sxs�JF�}q�urzb���sx�����V3S�N����y����1t�n�ayG��s��`Cʴχ�I�(�jY <m��SbO|�_FL�����^E��$W~WexOi2HQ�$ �!���!6~��4`V���a�n����P4G�<�	"qBA�V$7�1dk���6�섈���&B����)ם���4$w����m�TU}�F@�Š��<C˚.r�!Ֆ����6@gE�xիLVn(Q(T1εr�rb��V_Q�yq��ɳ��G�g(�*�	#���f~<c!Y�c19����s�x(��MQ܆���@g{�7(:6������i�d�0����u�W�Sg�ݘ
U�e�f�?T��z��[=���=�>;���
��oX�� ��u*�R�?g�A�㖣z+�17��/N�]lN���F�tmo����Pw�b�bJV"tp)��� �Lu��-��{����E�'ߖAO��I�>x�&����k&�Dd�(	�~�q�ę"��2�U��/���P�"�v�����NY���Jemq<�-Ac^��o � �
�;e��&�J��r�)�p�1/��,M���hٳ��_���^#'"����|�lJ[d�h>�`h�%V�j.Dӷ������bB���ƞq�}��ㆪjCp��0U�a�Sen�cG�B[�������T���Xt�
�)&�g�Jw�s�0b�6�bY�K�F[PS����ǫ}-gL�O�v~����װ$�zwHt��(Q0c�#�KPO,��ۿ�\��L(62���	V��z�(l'&)+�'W�;��ɿ��܆o#ɓ#�,��i֕���}����i�@O��n�V�K�h�VE�O&-	���xJ�^NJ��jaY֐#��2v��}�G����o��Z��{�Qu�ʤ��̍�|A�ń����1��r=
��W|��J= ˖қߙ{vwtz�^�b�k5V�MNo�+n�o���ڒ!����L�l�*Bz�X�������`aHr����mP���\���$3�9p+xN`&!H4����mDGv�gz�ўq-�c�&�˗`�q��"��ĸ�G��=��]Q�x
�)�[Ђ��۰|ɿ�0	�oh���K�0jBA�ǜ���0���b��Sre��Q��d��'�jH},���9��ݭe���m��O�ߓ֞�% ��Kd����M=���klq��h�;ߘ~�j\�g7V��$?M�,Z�W`M]�4Z)�Br�9���a>�6®H�&*Ly�%/�!�.	�Ȳ��k ���]������tW蝇�{;OI������77b��.����l���Zf�O�k%͙�n��w���l����Kϯ���%�\t	E�jHo�)I�"07{K<s�I�o�\�����g�F�x���)���%�wy����s2����u��/������A���d��'�u�L���b�ޓsTb�I�|�D��_���R8*�sŢΊ��T���'Q��:�MT��DR���#�n�?��(�T���t�o�4�vO!9h�;;���M�mc�a	��ZhzӀI���6�y�+�A�?��^ð��(�`7�!C��$�'*R�NXZ�����W�cJF��(&9P���H���o���k�(·y���|%�ͱ��?�����S�!@H�B�4��� �h�3�0��7v�=9������n3���fe�����sucr*&�~ZO@�0�����~w�r|۬VA����?�������6��lZ���L?�������s�\L�8��}k��e7`�*��pޭ@�qtM�[e���,��N�d8V.���"2��栔�]i��@����V�iX�S�[w���Vf�#9������V����Ǻz.��r�xC�V�a㨚 4@�~S�}�鵚P��L��ƧMΗAay�"���^��KNA�4�9�4��\�=��t�:���q>l]�G�&̢譧;��t���".�V����'&�I�0q�$�U��p�T}}� 9�W�D���Ԣ(�`���L��c�f��ؐ.�r���Ѱ�nM9�� ��7X��Ni�����[͆�}����]��U� ���Z3�YM T�<�K�(�3��������z��M%`��N�y����e�c�^믌[p��</�����@@���l���������0Y��ml�y'�C4��|V�� 풦s���ٌ���A�
���N��|�'�s��TV	��FQC#y��+6��X�G�H&ɪ�D�W28ち���
����4^g6
]��XѦu�B� ��N;�M����M��D��<ob�9����o���?tKa��̷�O����,�	.�d5�QM�ֈ��!5�3H���� �,���̂�ť�h�@%|�wt���sa�_�H �k@]oX/��#�P���XaA��EJ*V4w���R������� 땜��H�d�";��9b�I�x�tm0��W�˪F��gd�D�M�S95��v�~�k�����\�*�;�ph�d��R��UG��%Ѥ6 "FUDު:EP�A���jU�ȸ���4������j�u�-V�1�1�¾�BPq�SK0��`���2�����k;o�Ư�ғ`����Է^o�/^���?���Jh�`
ԃO���?�2$0ͩtm��9���a�	��F!�2C���N�?����ʺ�����T£mA���1�y�����lκl�ɥ���0��X��*� �D�O�j "��d������� o� ��YSD�iZ����Û�Q0��ʝ
����d:�2�z4~��Ъ�#D�������8ãZ$	�`�B7���|M��%,���d(4cn�aS�]."�Ɓ�"��^����Ծ~;�пC��0�x�{��}�~��8�����e�ik�߇:�T�������+�ᘻ*�9��Lo���Yw���`�94�#nf=��POƓk��@���VI���U�h+s�qۇx��gy��n3�#f#�n	�ĵ8�+�':��޷�����z�m���-h��&�����he�)a�W�;:9�sUjNE�k ��Ў#'�?����M�2h_
�O9��(C�p� �£���$��v�A�� ���]�6���rZјA��;��Og��%ې���Wf�߭�����t�� ̢�u�����Ȳ�	S��>�7���ܖ�g����&o��_�-��*��䡎ЁyQ寒c����/ʣ��V��W�
'mC�%~�����շU�����]*�z3p&���ǽ�LvuD5	F��9�0+��zOj���ꆓ��}�7�������u��4�+����Ħ�	H�����7k�W�ٚL<h�`:�,�D��-��V��8i��;8E����_VD���+`.��8��G�sl���	�_31=<ܱ
`�w�=�f��	��^�$|��8�o�pەڵx�����a�҉w�|*�ż��&�����ۓR�p&� ��u��-�D!_�bd;��C���sԜ��ցB�9�g�:�p�B��a���'�T�5<��\c������#�e�F�zm��Y���zb�.�rH�k��(�%����ș4�����X��"�����U��g��������,`s�̭�����&p��$ew�$���	o�,��Iو�j.�=x��������lf27kF|�6X�x r�1��VJ��������b�3e��sHXrb��x��4#�����d���xP�r?˳GɄ3+��t����a��}=��-� ���ZYX��,;��q�uphuBS�Bbx#]9Q�=�{�)z�g�EKKD�_*�eQ�Q����0�c�4[2Oƴ��[�dUN)�U�{��*���*L�L�S�����WL�U�����'"�=t���==���@��o����b������� �jyv5�wǘ�au�.����P��+T�f	~��>`	@�(�4+�V+Wˮ�Igӏ�`U���v���`gm��gб������XMs�owm��gXu�o��e�0�:H��S� '6�%$G<��U�(.�f��{ld~0��x,(�V�%J`�s� Mk(O�� ��_���QЈ�C{��୓���dx�-�i�՚%�ְ�F?7��6p��HU�5���v�v-��$������AAW'�>U.���2��m�
��!����}u�Ѝs��,��w�}�������bwe � �-�	1��T0C���Z����X-�+�m��j����� �����L����nA-��8�n`xND#��5���e����B]\���k^�S�A�Z�O�z��U�?��5�%�XT��w%�b�rҲ=�!䶃	��fvl3�&�������X÷ME��-�����V���ȀpE�Q�V���j�yc8�x�}Ŗ�و��W�@*�r���]�ƻF����i2���G\øu�g
�Z�og'U���i����<8�0�p�a����	���5NA����R� ������<�ّ��n{�|�l�Ov{�6��㥛~c#={2��ΙU��D.C��v��8�F5��X/������q�m|D�Z��jߏڨ���4�Hn*��@�u�l�U��/�EJ�F.���4�G�{�шG^��p"'bb����uj�.8��)S.q��O$�7����K�^�y��;�B��V���(��;���b?8^�kJz4���碄��
�MW���Mi�x�a�9WX��$�`Y4���>Mwu0TQ{�� ���-1�g��m��qӃ�1���B��AJ�B�/��pFDf�">�b�tvh@�z����_BG �Az/�Y�ͭL��A����:گ%�E�X��\$6(`�q\�7K,�9�y���=/�t���6��ٛ��Q�E���i���'���Ŷ�o�$26�5*��r�2�B���I��<�Y�Dp5��A�(�\���E��X�_��jY����]������{g�*nd�Aeв�z�m�%޵o�nDP����f7>e ��F��yv�o���R;eC� }H�9�];��ї<��\��հF_lZO��� ����gO�m&��k/���Eu�?-� M���-Aw��c���t6)����o��0c%�É��)�/~�AS4��)W~�{Cp��H{$�9��^��%E���.ٵ�{IJ9�0�L֯2�.��6z��������$�ܶ���Yr����?�R4��\<pa�^]�c,�Kqc|���9����8�0}�0�N`4�e�}�2��Z���[K~����Ɵ��Iz�;�JA������%47�	];}�H��y/���2�gn��FW�����4*F��vsm֞��f�t��KA��\�y�_q_��!�ʬ��B��~fa6�JB1W�df~���Rbp9ԛ[���_f��⿋-���/�h�;жL���{�i�5��^��0Y;�u�9'�,��s��4�3
H�gM/��v��)U
�s������V�0��^����� NkLޜ-��{e��qGi�?��,�+��q:9��$})x٫����1�(p4��2;�l���l�E������/�Rm�wJRrQ�*1��v��B���A ���Mz5?i!�&�w�-�V�7�|ˁ�Y?�bQ��(����-�o�x����ې��}�M�mH2�P��9��E4�pw^r�
�����>�6fs�a���Dj��uQcPY�I*�[����3s�Npxcu�ÂA��/�5p��7����6�<�͈|�9�c.�k��`�	iX쎓��w��U�$
K�O�M�f���L��pK�'���юʡ;:�<zc�籔��{N�HHvJ��):��H���j
�vU	����lߌ \�{�s�'������O-�{��ը2N�ḛV,�w��@5���HO�.��L<�H"M���>����p-Í7��%����ϳ�sa}�d�[/��k�K:�����2����s����o�'�30� ��m?Ϊ!0�О���Ԧ��=�$�����*�_:��J��� �q����N�:s�X��2m�g���o���_M{��s	΅n�
�k�8�~h'^7�m颸��?�������v�R��S�]跫�&�e$�D�
C�-�c��{$��>��&����z���Y�i@mx��G��1�js�<�W4ũzV]X�6����|���3a|�m�� ���m��@��Í)	�_���h�YB�"o�vA��*Ԧn�E a!�8���[��t6� XZq���S��fZ�3[�l�>V(>�f���!kK���=Ԡ@P����8��ne�p��C7�L�v�t@g�b��P�NNT�1��NXI )��	��
�={=�p���3*��w�i�U�fd���2��j.�˹߈Q�ߚ�O/�V��=-g����!���C"]X�R�s2�k������Vd����|/z?��#]_��e�Ix�d$�T���E��5a�H�{-E$��L�M_o�U����E�
Zq��!/B
E~Z�pb��+�G�
q���aH�S{L,?a��cNf�=������|޵��6L:L�d~U=��C�M� ��e�'���qap�+~*Vae	d�N�^�i�Ž�x-C_�$���pI�Fi�<$�)C�ғ�	�}|�����Ҿۘ�I����''{my�%�������8jR�����A��r
�<U��nj�:���@'<S���b8'u��NFGY�MD�������N[u,V����u6K,�1��CH?�ip-!���q�tw]��©�C���8�.*!���U��Jxʴ7,��yEVR�,��$gp�X���;f��n���Kr��h�?���)8��~�N��86,���z	���`��������cP]�a���Q�jxu�n�z�	x�-}_-)Ѱ�_z�|=8�/ �m�e�%=5��6��Mp�Ft��C�/�k��Oc����9M �Wu�-xKI*8Wʁ!i6���
�[�J�q��h�G�������9����"AT �uF�։��Z�%ݓ�k^����8ҳ��i��,�S�Ϟ���{�H�]rM$��X/��NX}9Im�K�og�?��
���t�?��MeϨ�Dw>,!5G��k3�%�ȇ$Y�}��!@U+0�� ��֪6���Q��LM�FESY�!r���͗#D�O��Ql�EB�
��i
_��˟��Dw���hi�Kb��I��k2�=N'jv�a`[N�KT6�z܊g���l�:�ir�:$3�^j��?c���]P���ԑ�Nw��V��8����f�g�W��x_�<�ēB�����& yy�G�byM��혇���b/�<?1u�O�n!1��O�z5�rj�_�)�ǜ�Ƙ�`f%tUDL���D�T�o�SD��{����� �z���Έ��b|�����u��-�e\�X���1��i9�a{��^BY?�T��y��,�E�C]v��7�Nջ���+�{��hFf8��So�&G�_n�v�c�`ek7!�U�Z&-R�+d06�Rs7^��}��d��U��$�%�z��dR�h N��R��Xਚ}�	>kL|(h5n7!�K�9G{���4����|�#�kx�}���o��IC����=��d$�x���!w����d6D�$�4�0ǝ,D�\�����U̠��:!}UㅿS����z�huk*F+VCc����G�c�q�J�����r$�Vt/���{�^�\,�����)1�=���>��(��&6�m�ix���}�=�E\����w��֓Q�th��D��D����zd�k6�*e����ϸ�oW쫥�M ��B��/�t%t�{��\v1�q�wo=��ޔvFG��[m�h+�;���od��Υ(���AE���-�n�=��+���/���:�h?�JE�>>��b�G'������?��p�,`8��e����Zq8Aw޹2���s/J 
����hzy��ZJ�&<Ŀ��%՜������Xx����q@1 /��S��C�1-��'a���t0^BH|���%� ,�#]��������DϧR�-�?]��YD����5Y@��ڥ�׻���i~˂��z����ա2�s��(���/.����
P<���~Դ.^'��z�g�TC
1%B�6_.���̘D�I/���(��>��{0��;�$R�u���ƣV\*��;b;]�_τX�z�ʧ�h�2�r5�sζ��}P�/\]BW�^э���v�G޳�|��j����V�ݿ��-�	��
�qO�-չ�ٟ[F�03���+�cPS�@>oV��^�E���A�� ��h�@�Q�����-������T���o���3����4�;�����9�Mt��?)'tΦ�0�8�.f�H��kU^E��Ӱ����O@��DU24QH=�ߜ<���]=Gq>|���q��s��
��pL�J\����r���g[A��ļ�B�rc>Xv"BPƌ�u2x�,�-vv͓��mO_ʀ�P�E4�Rz~+�P�๵X�{:B�TA-V�i4q/���K�#{�5(̕v�4�"��:�zX��K����P����V���ƒ�o�d_t�C@����b�O�i�.�����SP���R(س��$!�U���A�v3=�w�p=[Xڹ��T��3���w@Y�û:����>���~��O�&��Ͱ`74�����NVؤ3H�q9�w �:U�"�y�3�H�Q��~�_�T�U*	��Cէ侣2��}4�z%!҉�L�Yڈ���[�MQJ�9?é�7@8Z��	{ ��'�x���:1�j���:j��e���9W,��*k������s�_��;uJ��g͇$�?�qf�G9�[����8=a�U�/�Z���?��Z�o���<w�k|�T�&�X�ZRw���_F�n�z.�w��J��� �H��'�Ò��0왝K����F�=��s�$v��ه���7�:�i�Ns��kq��S�ˏ��jx�5K��p���ؗ5��7���Z9,|�sv������1�7U����壄�~�ĸr�f�'1�w^bO^q́���b��O�9`A��U<��lz����̠��q��C�-TP��D>D�Yc�R�i���,O�34)�u^��ou����:��ߎ!�hH;���j[�'h�bﴽ��r)��2�u�wO�,02.(�I���L�� l}�1[Jǽ'_O��M-��e;�����Q���ne_���W�Yy��+�X�+�~F�-�����$�}>ټ�n7j����u��VY|*���qf��N 9�/ �1�g,�GrqP�C�<���(%�C!{�ǒ Hi]v?f��� �S�����!�f�%q���U���#[�$+�i����h� �	5�뾢Q�/s��6G�J�0җ��smHԲ��Bn��s�'h��F�I�E��R�����Lth�r�Y8� ��D��V���]�d�jLPk���Y�1�ܮfXI�n�K��9�S��G��Y��L�=Nx5�-�;�d\��	`�G+�9䗞��o��a�fOauy����4
Um/��[b%�����ᨖl�!\V�j�����w���ްW�����K8�6�~�~��Bp�y��MUyyV ;#�n׳�ɖg��ܯ����G�[��&�E�f
w^��RX-3�^�q��6bE],B�>�-��%���OE�1/�1ªD��X)}a_W�'��!�4�*d�#Ѹ_�x����:���=!���bӈ��\���;5���
DGj��ɨ���c���1N;>#e�wPV8�+ξ����ۻ�C���v3���	^*/���.G�b�I�����˦	S �iJ�%H��a���t\�_�J'���12q��1�(����Z3�.��_WQ�]
QU��'�xؚ�n&��򶋏E\۸���q$�G�Sy:s4ҏ������V,��e�
J�P��x��-� �$+On�Ųm��م������*/�9�%�3	����`���l��Mg��_�W�Ky�})�����|���G_�)c��-��WY_Ϻ;��w8#d���Eñ�F!'�n`%�;H�yb*D;N���37����-ڸ��2G��$~�����IV�����\'PT*������y� ��ܰ��$���1)v�*������y��GJ��1�J�-~�y/42� Y�_�Ed�dz��il��OO��#S�Z��y(����c���l��DUry�C�������0���]_��fm�YL�dw��� >`<�&
�-�DՏb���>l�q蘆��qrP�kH��~�j�60(������,B����L$�Ao�@��4y�K 0�'���vz���A��~�yN�p���N@h�lOS!#R��\JlW��]�f{��+4_p���3�Z4'����ylq����hv}azn�]�́����3xZ.0��9���#�k�c��e��A�^9,&�����A�f�U���صK�~<B3��n���#���xM o��|ކ�Tql��d�)�/(����혗�O��W��w��eIpA
\ؽ�1Q#�3+�<~!��ܐ�K\��8�Wٛ�S�؋{0j;^�?�C��4����6YR:�W���1O����l�s�g���L�E�dCS&\.ڢǮ�Y��1Zr|�UL�;8�E�u�2D��o���m�����@E/���{�`�7�`ﭲ	� 9�T�e	x�.��Y�T�_�-��ɽ��Ss�&��4	V��!�a�x`#��ƥ�YT�95�k�f�)AU��(`�����c��yv�s��ǁ�ޡ��?�6��@W���[�i�"�O�ٯ�!QX��lZ�, �2ɑ9�fQ;��� ���_�4�^�8K�?I?74;_���$sr`y)+��yP�Y���@��	`b\�Ȯ����iM���swK�ʹ�TO3�NV�f����֤����w�d�j�b��"�3�(�_���F7�b��H�/�Ԛ�J�~�;��MD�ܚ�C�)��2���NW����F�.���:��n{�2�@�zgx�C����*3�PD41G�켸w���h�o����(���LO��'����$���w�*��fM����-X�ɏ��X�"��+ŵl�r�Ǭ|�_��\�@_�0��o�(~~Ł�B?2�p-z���j�2d��-���Q�$x��ew�	s�e�N�f7Gfl��d����}���!S�Æ�xT�S}���ô��X�b��kX��qDD�K��4�˻@����<����}�ߌ����ޜqZ�������3�E'Ir���51��(@B0�k�6�G�HA��-DّaQ�,{i�(��M��8��?}<Ⱥ�I�(69�(Q�����Un8rE'�;�����^7�-��ȄbZb��'�׫\{?�Y��S"�0],�+���X��M�7u���;�������bd�Y^��m�մ�\�������u�������e�Ѵ�����]9/����/��0V�,t�m��ˡ�� ��1�,s���R*��~�&_�-�?�Y=�[���"c�_[V�_��Ҿn㧼V�X#��1)���8vp&��B�^iXt���S?�K?����i�E�
F�'�K�!z^�Ύ[�_�%>�4>�aQ��;fSU��O���$[F��{%O��uj����MX7�D+�.�uϝ4�im6u���0N��h�뺩���2.�p��f�����
������m���q��=I7:��%|`?س�K��� S�6x���P�vs��ԥ���BƩV��#E�t�2���5e����]�x��������76�z�E��$���-Ex��I�wQ���%[]}6*�������_6�&̰�k�ySa��iO�֯r����z���,��l���~����@���}�Pdf�����.0��͹f7+��i�Y3rLQ 1R��k�4�-�G�~�����VS�bo���lX��.-\�D3�C�Ɍ�@��/�ޒ�|cX���2�;J\����]�`�u!��lW�T��>y���\& �D����NLަ��64ɧN������[מ��C��[�2{�SQ"Zt�����L���1kg��������|&#��蹲�ɻ���>�\3f|�[�P�K�;
���Z)<�C"nv\K�E�j[A�ɾ�:�m�p(����͝b���N}B�d��r-O��ǼA�ރك__X�5$��߲}0 ���bݿu�:�^���= v슅������ٿ|C�fpa�=?�����H��ٯ�����H+'��J!��$�>��d������a���4h�}&��i@��V;��h�4�x���&ç;�Zն�7�7F���Ծ��Z%�gʇ�jY5sX�$�DA��b�)�*�$]�4N9qn�o����ӬI�cϷ_��ϚR�
y����U|O���lN��Н�V�F�퉻Pp�c!��̀)>�!�^%�$6���N�LG��.� ���S@��.:�\�#eP�+a�&�L��e��XE<2^{[�� �����]��l���i�քZ�{
�^��������Ԛ�`���h6�LN��u�QO�J�Aj�e��Q;��櫳j�Q@��RŖ�HF������A˶�^�6�ʠ�BB����7�]$�"�@M`B�(���u���b���2�V�Tʭ��R�֠�70��C���)�P�+1�O��i������y�+�LW�`0M�M��h�]W5{:���M苰߉�'}͑u��U��&����g�.�Rd���M7��a'!-�þ`m�k3��x-Ss��<��_Hx����\ː!�F�c�+����D������+6�tZ���,��(�"w|#�8f�&��F�`�×�(�|�NԘ�U�UU�������"k8�� ��a��V����K�<�&*���辘:�����Q����"�(� �{M�*n&���A�_&'0����#__�hlh�sg�g�vbo�1B�Hp�Hc��/���`6^�@�'UuO�L�z�n�y��]zL�E���j��KԒ��%`����{��2~sVl�g�L.�ݳ�\�1�ʿ X��Z��i:$��榑�C_�VP2 ��V�=;�o��ǉݦR7bl�]�	zL��ѽ6�zX��A�K��**� ���鈑ɵ�Ǽ�I<��0��i�ܫ�k��}��n��rE�A����ȁ�!r2������ة�t�������)	�V�����o� 8x��>�ǿ������{׵,JV|����Z_�'��V�"&3q��n�����I�P��	0�[w��'��`U�kB@�<��;{UE`���A����?���9\��qw��aW���|U�t��eycb
Eu��\��+�qg�6Z
��wPIn+|-3����g}�Z�I��p>M0{�����S��{��D �ʻlro���Y7��&���L܏.ң.<�!�q����(���woq�Z�%���o����򎰏�ݷ�+ �u�zى�R�Av��#mD����U�ki,m�s}���U��G��&*G��!���TwZK������
0��?k��_'x�tyn~2���94i��8o��w�E�0�X�ʵ;�lLҴ* 8ѥ�UlhS�D?��d'
z;kft(�Y|x�Dk]���z���q.潭��@�W_�;�My�L���Sͭ,��V4t1d�w��6䣮���ާA��g
�߽6��l��\R�Ս�6%9�{<����7�<h�qŒH�@x�ѿh.�G�c&��[�e/��B�5t)���ڝ�g������;Y����y9��DE���`3Ĳ��'�"�����]A���
}>=�3�q�I;F��:�?0�+��C��C)��_lR�V6�?�Ś����p��H����A:��6H3!)�Z��x%RS�T����:8���3�ks*�̭V'3m�P�N[m� g���������JA�Ј%VKH�%Οw`���,L ��GW4��dܥ䡂'���7i��\Y\�����¾�2�x�����eBֿ֟Yے஋mm��B4�*�GڑGr�y�K�k��օ��X�Q`�qٿ����KUƒf��h]�	���ώx�����,�~c��x~��;���(��Y���Sś~&��P'q�y)������~�� #K������.�S^<��c�aR��P{̎��`ի���=5��Go�z�E&kQ��%�p��c�3{.����}�I!L5L-20y�Q� ��.�7TE��X�K<��C�J*���#�6l�@,Ҝڝ�Y���EN��KR&��\G�-w1@��Ae���Ms8�>b���q�Je�7���L<;��{�\�)/P��c��5�X��G`�� �|�?�E,��I�1���h8�.�P ���Z�X��g�*�=O�p����Zɒ���)�*��b̨=�ӵ'��`M�2���؝�s�-n�tY�_AV���UQ �*��Xh��?�S�v�(|<Z�� d�뚐5.�'���)��E-��W[��
�2E
�I#�S�z�7Wi�L��s��ۏI.&<x�l��ߢU^�^>Ț��M���~2I<��ͯ('�qj��5��l������'����/nD>P�Bzbuj �J�O¦��$r�
\��g��9'�[�t�j�֮���ur�m��3.u�O�F�I�G��R;��5r6�$g@<5x�𢅴Ṕ��T$f�����BY	ކ�� �[�D�E��]�C�d=��\k�o�#���'��-4r۫A���w�}������O�oz�.ḻ��8[�$})|ɫ�>��Mj���:�, ;-�I����p�e��G�=�ר�?>0N^l�;�MGOHC$g�F2�.R�������r�;�Fn�%EK�N�JK"jKY������w�`�?�h���,��������E�TN�m�#`�b�(�>
���☤M5��S!*�%��񷤿��~��E8����c����mk�nՍ��{𞙷G-�2Eّ�N����њ��U���g�����'{�ڨ�����]�o,r�լ����N���,"���f<�ZVm*寍\��"�*��k��Ctgc�(������4데���ȏz���r'Tp�DV��W(�]R�3�nÕ�F��e����O.k@RY<���z�E�=Jd�%�����
^�l�V{7����M�Fq&��!x?�Y�J����k'�$Q������ͨ��7U[�Ŧ��y��/�T~�I�'����+O�H�1k�8A��F<�I$>W/oU:�气����O�y�0@�J�}/��:�g%立R]ER���y֔G9�]z�jν+�������M3.I�.=7+��uW#܍-�ЁM��Ib�V����z��������nBg���(�g,O�hf.|
P,�5�N�X$^s�y1���RL���C������ነV��}d�#�_� FP��#��m�FL5��j��iʾ��	v�ij����M����]��'tQ�O#*;�6��e�e|�@`�ʿ��JX(��Jy|��3Ms���l�ڙ��h�*qO�&��u�A�)]<�;`����Y�.�o��dC@�T�#�B>K�`OB~�d��ac5�@�H��[9@C�$��,�y��M��������o����m�r�q��&���+\.��B�9��l��(Hmz������2�<.yM�I��;hۆ��@P�n����p��e���`~[BL ���q�1�O�{�
7(�z��i�v�n��C�DV}w��f$���@{���Ao�@�����D�q�1��	P8+E1F���Ҵ��3	U���ܗR,�����N殾۾��(5�T�C��M�!ћq )@v[��`�l�m�Μ�f<��獥��N7	M��Y&��"���9.�X]/����.QK��+o���3�w�](�<�v]2�DI�Y��"X4%?�wduz��[��x��}��no!N�̗�(_C�˧�2��Xn�Up�[{�
ub���%�;�jv�d�gf�	D�#�0e�9u/m墆�+�O��aHY�٣�3C��]|x�G]��u�ď��9dwO/@c��,g����d�SGɿ����'��D��l9�/�(b�Z�62�\�Do�1��f���`AviR�Bl"?. t�����?���J":��( ��B���ѰR�ݬX��X�j�0�%��ɞ�qJ�T�������ޱh,S^<s����	�c־ƻ�'����ȫ�e�����+�O�$�ɾ�JIq9�<��K�+d�9�h�1���}Z�ּm"~:o��O�)��R���[��d����7�ŚxS�509q����߷j�����e`dՖ��[�Y4���JOU�IȽ��~D�2H�ۂ[�'%@���֬��~�0+4y���yc��!*���,#>GK+���j�O�@���x�Wz�F�����q�H�X���ݝk�HW���]��x�f���Dz�ż�_C��Q��74��_���b�H��i�[��J"G���Q�N��9
R�޼��#"8���V�L�`�	�k�
;���t�N_�;���ѱ�_Y������{W�2-��R����A���
�#������B@g��7��P�?K��b|X_�Ũ t�BSTB��Z�y)�?.��5�ޠH]�������V���n��ҭ/������ Wq�8�	�ȶ�������1�FI.���'s°�O#fH�~y��<rw:���ОVD����q�R'K o�����l��taѧꨕ���\a��AWC�۵��!e*Q��ޅMO��:�z�θ�>��e�K,��)�h/��(lIx�����^p��!��զ��ץ�t��(��?�S��)ܻDs����]�k���˟�/�k����)d� K�h�ax���a�I�5�sz	7�vѾ*#����0*�L$A��g�X��^Z��`d�(;�.����0�>��9xo��^>���7�g <��5zg�������?���:L�$�e4�;�	�������<p��`�%>۹g���~��K2���!'֠BHkΌ��^��Y��y%D��_�E�������15�s7+����˥�Hg��ͻ���L+�h�D�.�7��2[�fl|��`�������D��ȧu�]UXr���,��5 v�)��"L_���_c3��֜��<A@��M�c�Ը���֡���Ff1l-���B ��q��zG��Ϳ�̌P�m{]E�;}��S�R�(��*��WB1�{��i^O��= bٞ c83���W�	�ؕ����i�OIj�oQ[��$���hrΨ�i�j��N������SL���̒��,:�/��@��۸"���E���	f�B|�Ck�c"��\y:��Sq���#w��V@��$���V\��ۭ"��ҿ�R���������D�hl%�dXx��A�g��y#��L�b����3
ʗ����D���6�G�D�:2�#h![��7j�%i8[��5���Ӝ������P^R�/�<O��L)�f_j�� Q�6�ns�d��Q]]��[g��쉫j��G��G3��m�P��k����qч )��BsDya8��ZRS}�ev#ȼ-���X�!3[I��*���j�@C&M6���I��T�+�i߷��o0�vbp�Eil{
E��\Z~��E���SFԃQ�}G���^q!�-����k�m�μW
�����H	U����LdqX''���yr'.�B�s��7����-+ċ�DX�S�|)i�I��"��g���h���X�pI�GqFt�OLV�Q�P8��@�R��������f�kH�ՙ��P5{aM�SXes�$Pg���V8_���^~v-s�i}������aP3U=�
4y�& �Ge'�p�'�s���ϱ�YA�
��\�&�_�")^�oxe�Pi�E��V�Z��5�r���S��Ӥ�#z��~w�HõO�I �nn�e!�s-�]�V�Y������l��Á���o"��k{P�:��k�gg	Z\l�m�һ�᱌�%�<��ZwIY.m���N_�VI��oT�t���T�xB��Aط��=��pr�Zkĕ�Y�"$�
Y#�u�`k^O2n� ~t*o9���Vm��	�P�t�a����s�lB�TO��-�aj� K�"�Q;$�,��Q@-���*G;|��׵�`�%��X���nW���������Q́ʡm>�x[@���/�kO�i���*l�?~��q@'�dӸ�%�����1ϻ��`C'��՘b�Hj�`_?1S�^:d��P��7�a�YC����\�zug�J�A�$���hI�U���''Y�d��(L$���@l:o�L�s�2����gkB��Z��}(~`����۹_ּRO��g�?��u��pH��-`�.
�6`�3� ������X���Y��M�c~�{~I����n������]�N���72%v��5.�ɤ��(L��q���#'�q�+�Q��a��hƫ������;5��ak��&�0�?�'�>�L7�e��N��y&dq`'T���c��be[mʐ��e�$����;N�L2��{�:M�\;�4:�W������W���A������O�" ���׀��Rm]�qCҴ��.�Zsq�n�?��r[���6D�� � [m�������ȼ(����x?�B��`� ?-D���-����/�xu�c��tG��ib�v�_<@*��y��K�a�^�:���I��Q�7����\���	��0h�$�1��n�O#k{��]������_9���1�6�f��#�6V������Í���ܬV������ ��2l��߻X��)��N:��00�凾���������/�n��K�;)�R��sk�����9̜�N��{w/T�^�K��&=�D���2Z?�޺'Si<�j�;{5����#�v�6C�i��3����!�;s�9�1�t?�Z�;�I�8w���,�����s��3h�ם�:pXKa������āxҏp��S_C9�  ����Z��ֵ�L�Q��S���1T�۷�1@v3������R��>0Q&�(�4��y���b�Ԁߨ��\$lnq���i�D��Z/�_��<].<�8ҥs5�Hȶ1�%�@���Wt1&@UR>qN(���dV�B;��i(�u�m����X��P�i�������G����x�:�J�puOv:��0�I�K�|�>�X1O����Jp��rR�ƿÝ<ܕS� v7c�)�,�UL��c��b����:ȥ��y��N*R��>s����ڊ{<a(��~رY/��L��@�B38\p��5�%�ڨ$z��8㑗���6%k�����Jz']�o�������E�3̙��q�o�#���c��z��q2��'$���e{�c�:x5�V���� �T�2�]s��N]1���t��"+��If���Aᠽ�.S������O�x�����`.?<i�ז��{�i�In-�k��I�o��J���@�"�#tW���P �� �� �h����۫��4.�z~uZ��N�w��Jo�S����)�ue� ���2e�5��0`1�*���)ѝ�g�a�OT��Ϲ�E��8җ�OF����������71�!6
��4|��B24�D�`]�IK�%�E@I��J�ԙbK�< ����A��H���:�W���*^��f�Q�[?d�,��>����N����d{���Q�@&Y�Ϸ;I8(��u2�)�u�p�+�0�?64�R��c�}�k#�@$�Rp���u�L{0L�򓁒�o��c�Bu�K<��O�a���j�s�9��Q)Ff��jqA����52��j}\�z+pd$�av�¯���
m{S�5#�mU^�a�n�E��
̙_ě��\�S�Q!/َ���=�;#�gh��HR�h��������B�(��1v�YL�	��Hd�Ce�f ��s[�bK�{��o��[}�
�xO��Q�	�?���>�/��H�^�M��&���0\=�><�Ǭw���m�!k�|%��]
e�p��y��c9N���E��'JeBv"�-�Z!�Q�p[x[�$�,瀢ۍ��W��ǅ�w
�\�+)K�Vc�P$�o�;r�$�oC��|�QkE~z�B��k��+v8߀&�m��-��B�15�*.���a�L�"�J���"L��䇣˞j�c7�'&���0��ն5�P�t+Q�X�V3���?�3GYQp�h(��ֿlO�d���4()ZL��ZHjA��:Ny�?����EL��	Y���7q���~��U�+�GkO�� ����w"�0Q����4T�G�Q��|:F۹�9f��͘��B�t��5*&*90�}d�d**�W����K��R�����0fo����#ٍkگ�Uv�y#����,Wh�n%&�{�^_b謮��2Jb5�jݚ�Kfƛu��~���璱��"Е��=�0>��t�6&7|����wm9T~�f�L�ڸ�U�/�V��������������O\�1rX��;�w���xXS����7O�4����U
�sN��Õ��߾]��t�4}���Qbϱ����ޒ�Ҋ�۫lX��� �Ha'H� 5��>a*�E��@���2d��8ö͠�V�x$c Of]�6����s���7�H������N<~�O'�5����e��Δ�9�~��J�m��^�$d���}���	��ީ��`X�-{�����V׌�Ƥ��rZW�C��,1~X��=B����GAU4�=��� �cKz�z�a�QC�/��F�+j�Ju�qk��'�G�H�������ۼ�H��Ìlh
r��U����{č������6.��m��Ѯ��ۃ����k��]��;4~K��G��ko��Y���
kF����FF��mM��)����P��n>m?&�D<�����'1��Ν|6��h��Z�hN�1�֒U���
�h��:�P^8�қ�Q��ҡ����b�����߾�@������� M��)��.2+�����|F��<'$��__8RЌ�&ș&�#���aڋr��U�.���Z��+ �J�ko��(q��;mc#yX:��*��Me���hłK�fTa�	\�9�mi�Ex�TW�(M����S<��{H�[P�?�g	`�5J�i��j0`ɣ��Y���&x٥I˟�s��f���z��f���If��6����¾n~�Z�xp��Fn��|��@��v�!㍞f�6f�.sh���P��@��� e��Qi�n/�	�F\��<g�k�q����[�p��� S�T�S��(�����W�3-�D���Z�Ӛ��Iծ=�1JR�۝�ӁzJт�DX'���E���|����t�z�pK?�YA��1�856��f����k�O�NK�yr���%v�g��<-Ado�e���W�:͙R�4DƘ'�ޞ�z�tp_�!�l-Ֆq!%�2B3�upᢅ�����9|vn� ���q�D2�<r����ni��^����M�x�1��7��;U��7E6�;�B>�c�oD��n�<����(W@B���"׷a3w��G�v���4+"��s�KGo,rk�)l�<�7�h[��A�|�f��w���>�z�80ntI�^ޡ���X4�u6+�����^��NT��q�N]Q�����F��R�@naڟ�����Dڨ�y���Z���e0o�@�7���K��(RObb$s Y �8�8��7�vX%��
;Q�yZ1�+�Ll�=�\h��0j4�e�ɂ�u��-0�q�sR!'R��?D�����MQ �w����QB')ϴ�X���[2K)�f��=��J�]��uE���i��S��Eݼ7�²:��V�@$�S����ٙz'��"���&^*y��g}��E����X�c���Z�9z�8j�2V��q���ۘ�&�'�� ��=�D��1{�0$�A��l��:s�����ʦ)�h�8�>>O�}P�Z��%�O��đr:����~K���#�KU5�F���طu�i����f�)��9�������ܖ_�.O�T�
q��d���D���o���i&k�U��Q�	�s�L�@YW$�(��Ա����"
Z��P�xSw�gQo�S���^*���;;��Qo�����
8s�!�$4Y^'��u���S�؄av� H֊��*���������H!�b���D�`�%��F��	:P$�pA'��Yyu ���Y>�%���5u�h̗#s�fA��I�6mzjk�Cp���,���)�ջ]!��.ю��h�mǡ2��w���i���|3Ku�\#�1��xK�`x�(X�ݘ�v�l�5��>��v0��؂Oe��"18%�Z�Hl��
�\E�9
���Ї~�>O�9��&���:�u*RF��sS�11id-2q	\'�����^�hϭ]�*v� E�ۥF}���\Z��l�Y4<F��+��0��*�]���0u��}~��~�9�R��M��h1sTÆ�p��L7)�%� �b̚��p����������:�8ٮ���΀{zv��@G���v�2�蹴���ᢕ�M�0�1�����!Uh�j8󃺕9B��[������Z�y���p~�����N�U�w����3�myz�-��L��4���;`o)�5������q��$}�Mn;Ic��_�
�O��1��UgQr���+��(;�R+�nJ�&>[)N&�ŕ���R��&RB�mb/�[�-���vo��(�>A��R~��=�1��t���!�.Gd�����fi�#���'�y�9C��_����*t��#���@<�&¸�8��JvR,�8~t�[�ׅ3��f�y��j,���D{wQ9�����Z�"K}��8�*H7egTxI�}'V����\��:J0M������څ�=&Oɗ�|7���e�V�<طK)}�p�|�Dn0�����o�2 �8���S�nM4�v�xVp��iKC�mww�d�&CB��Cv������������H�=ä	����ZY�'���*>���T�������Hf���+��L�c٥0d���7�@&��{L�8�~��Q@*�3��h"����~	�*��Ho
ֻMl ������@���eGQ��⯚<���%I�i�WO!�>[n|H�.A�� +e{��}ܚ{���O)@j�A�q��J�f�=� ͺ��>GB6
ꡓ��UW~kK֘�,��4��)�kw�TGW�)�',yĭpM�@��	��@m�K���Sx������Ц�:�>�Nk�p��f[eS��8�������.a��8�P8TL���'d�W�R�m��C%�#46%�>��(���Rþ�6i(~`^|����{^֦ ��kJ�[��Ǎu�;O�y�d2~8��_�D��l���)�P����xm��|�eY75p�ޙŘ�C8)q2w� �����w8bΥ����������v������p��0��+�>C��`����m��)�Z�n*�^{���5$��k�{^��.M"}"��!���Mr��j�BMK�%ڻ�^Y8�}�&u���?�sSI��5�p@z̈́Z�A�MJ�f�rt+-�]����[9**7$G߮�^���g�#@�L0|����hpW0��Z-�vB&�u�O���.pI�����x�ђ��M��+	l��+�'�k�)5�B����]O:/�g�� ������e}��
V[w@Gj�;�ъ����.��h*{�,6$ф����w6�8���&�뒇 ��>^Z�8wh@@!�h��݇&6��[e]h�Kj��e(\@�{�s4�A���P��g��P�5B��cϿD��������`�z���t�k]��EJ4�	�8�S0��!K�=B�}#Pd;����Hm8$Q��v�8�s���+{K��/�#��Z�w�ғִ�����'ES�Uy�p��O���������9�^��9|A%�g���-Ʌ-*z<6|��w���@��5�R�?�����UM���w���h�C�ڰ�R_�q���Ÿ��Vnd\J�i㿬&����{�����7ׅv���HI�%P@һ���'�����DXQ�XX��Q��>��"���� �F��"�����z�'�}+,z0n�J��w3����XԼ����\ww��@��H�Ķ!Ŧ��&Gyit�QsX�i�HPTεJc�ߡ: ٶC�5H�J���m�� �u��7)�+�Ku5�����@G�K�+�eW�Mپ3C�${���2��%�^��-�M��_c���5�f�U�"&��GV��HE�`�ȹ�(�Uc�U��с鳧ݶۈ�M�;�������҂�0UL�ޒ5�ڿL-=n�-���fuM_���c�VK{�Z3V̫�&]ΰ5�)`/j��Xs�>7C*����`���ɵ����ų����_���Ia<y�)�yZ�V�-�4��N�Bj�g����;�pD09�2:HY'8�D(h;����H���>F�am^f>�嚔�1z�bpA�޸�7)єLQ+>��4�.I�6((/����S���>��tXٟk���*0q2ɐy�}��qR8���Y�G@��;����P��V�q��K���5�m�Y	����o`U?MZ�����)䑧Iq�.��:���42�40#1�	p8���d�*��u�w�����\f�"p�ܑ|)�v*�f1'!	�{1�*�4B���ژ��X�(�"���%�� �z|m��e�=��I&Z��t%�2��N�c������JYe�0�
V5�ł�: �e�������M�ͭi��2IA�"���"b���v� f�~��	Vc�Q|�{�f�?����k��P��~m[iL(�X5�Ԩ&*�;��{nD|ɺ�a�ƻ����w�h�[-���Kт��4�H<B�)HT[G��� GY�
�F��k���-��@ģj4(�'�yb�"%EW�x�������]�������|�����h��͘@ͭ/�yy[q�G��A�
�<(9�uL+�y�M,ߩ٘Dj�>�����������+�0R�>׺�56������P�riF�����Ar���	�\i9u`3Y��|1S���|n��n�3TuƲ<���P��é��;����'��˒���dD��?������9BZ�=���ZY��Bq�\��?�g3��33�=��C��G����{~(��Q��\� �z�/w�C����n�m������P;�S!�Ƹr���f�3&���t���c��� 9�_ �רPF�@�\���f^'���ʙE�VEn�8�e`��Xhj�D�`~���<yl5_���8'�0�`���_����o��'%6��<,����Z� 6��P�wȅ��3���������WDyk���i��SУ�JD�1�vT���0�eb@����O�A}q:-����Zנ׍m�m�V�'�E���Ӝ%�L��T0�K%N���yH��4d�������^RW���,�C���D�ۼ�gC�Xj��>#ù���L�&�5��0v��L��ږ:�>8~���8!�ʛ�đx1۫C7,"���7m���u̘�I��g�N��P��|������S��$�:d�����5[��b.z���,OΧ�RB}�A�Y=�aq��5�FyD��@�3+Q����TI7ӄxT���U�
�ْb�:p���#��"#Y�\?��'��lT����C��@H��t�����EIY$�nP	,us��w70:�<�g�6Zw������$\�3O�%��CkC��?S�$欩����HAlA�7�v8Dx�,���ǐ])`R�8K�p���&1 �mj!-�ݙ���hY=Z�><|`����t/�K��.��(�&����A��Hz�Б�ǤO,�E���9Z��Iғ�f��
Ȫc�2P[�Ae!W7�t���.C��?��W�<[X9>�I�[���Ð>兀�ҽB G/�rɼ{'�|��h��7@s{A�Ara���x��kf�	x�4����a��G��o��+����4�'Vi��/��h���<���@g~�<+��s��`e	r O��Y���Ó���ɯ\ށ&�obk���me��҇�i{)M�w��40	#��8�g�9���^�?0���B�28i�^c�[���QX$=c]�;`��(�l��r&px�j��#�Q���4�c�莐0�$}�>����yRU����O�͑.�S1q��T�ƼlI���m�u|�h�".��<J���'=��|��P���qL;���3v\R�z"3\������I�i
������u���R�C%�Ֆ�������;��a�㽐�5�~3E�Y4x�(û>�̃Q��W{Ȗ�������(N��ywȶS�z��ʉdF���Ƀ]��]CYk�;_t��}G#�9b^ld�7�)=�7/���C��A��5��.�DE����0��Ts�D��?��Vr��Z*
Bߖ=��{WC�'��_�B�/W�j p��é4���̵ ��G���(�2��$���Ň�\^e��6쩕��eS?u[B�i�P)�Qщ�r���r���]��� �M>��r4Zq���y��[�V?/fֳe��	���)'�{d� {h��5qF�ƀ�H�
��fc:��*E�=J���J�E���Y�����4���^i����ԙ�O��4����h���"�+������f���l]_N��e����O�.TE]v@���P"�C��I�Ս�4�� ��)�=vup 7֙� q;J��w��I�$���ǼB8nF�\��.��T!2Z��p(�� Y����\C1��j���p?
9��f_��i��J�LAx+���6���_L��[k�"A������6­1m>T\�$�XΌ�x�ϙ
���=ŝ�H� A�-��+X�����%�ɚ`4 �C,�����4IEf��͆C	8���ۖ��Bm�e��"4�B����q��儑뫰���;97Q��3*f�n8hH|�kv/ݧ�Z�9��U�,\x�h4��-P.�r�K�hM
r����o+�������
���&��F��g'{S&�Q]Sڌ�Gg���6.r���{f)��:��Q��;�i�y��AYӓ�b�"�t8��� ^O5n&�Zڵ�:3�#�["D�����?-�s c�+��2�LvÃ�;ej�J�;��E��w&Ѿ���5a�!��;�.ړoAQ�62gf���+|�Ɠ��1�w���o�]��<��(=Sj��w|�O(��~�Y׫E 9*��������D����"��D�̶|ݦ(w����M�f㱨%�ܔ��^b��x�_�T�o�S�s�+��9
�kW��E�gM�-��&
	֪�g;� ��V��vд{�W1��V���>k*=�y�h?�s���d������Fɧ7�6���b�����5����tx�|J�<,�.Q�q�|�Ī��*G�"����:o~��^\G�c�q7�K���>Ϙ8k���P-7�o��vɠ�h��rPj
�˅��k���0� ��l!+���V;�₫��/0Y�5<�&���7'�|��I��1)Ӯ�vDjN)/n��(G1i�)4I�&� -���=��1���q��V�a�2�Ks���|��Yh�E�T�woz��ӛۙ�����)�,��1\&�'s�d��`�|	;���T� ��"=�܋Hj��Z��jy��Vi��;�5Ddz=���%�����ݥ������PF��*C���v/��ih��Ͱ)IX�-h�^
RC�,�d#��̢���R�R�zR����������Ƞ�K=p�7z!�#QAR�j�� /���~�p�t*�~� ��N���-@��$b�ʊ���,���9�
��m'a�L��~��[��HpѴ��3gMm�DTƦpj�>�ĸ���L�����]��&$�{�N.]>(3A�SC�����\̈́��s���n�������)#'���:��(���|D��}��B(�]m�;`Ê�i0`�z�?����p��I�C��.����7�E���*��{��Ֆ<K!aL&fI�!��Y�aT��F�<�Y�C��  ڵ��i�Y�� /Z���̻4�-�]*{<k}��E�j@ ��be�i,�Өz@Wǉ(��Jc
��c^̲��<�&٧�s ��d�>�l��'|�8}D�Y��{��)lH����SрN����w�Q�u^_�=�n�htH�jp�B��)��RPV���,�U/~�.�'�=�8�Х@V?�f��ٍ�����nK��w�Yߡc�;��{�a���@�-���C�{rfe�P���0&\9�'��?ğK-�P4��x}��%�k�+vj��"��<�h7C;e��T����-t{ò!����T�6+s�I���\�����H�u�"~�^څf�l��[R�PGY�E\I��m�h��lAT��Q��@zU��X�MJհ��Fhj?5�GL�H�;��*�b���^ߑ�� i3��[��V��2ݻ�(��[���M��U�2�w��?=�SYV��'��9��Z��L������"ƽ�7H�i�M��� rA?�����%��F\�sqzǡ������U���a5PlJ� ��Ev 3>����s����N��"/j�GǦ�wZ���:*c>p���=�S���,�1��/  �E�Pp�l��<�?%`���q+S��R���D����#cepO��}�k(E����o���W�ə`?'�!r1I��T����W�T�� ��qE`�� ��^t;�� ��]BH�û��^Y<�r���d��w+�c��m���}��v�c�zh`�ۭ��f�(O2Zt�����e�{I�Hl�c�z<K��F{OJ0�j��7HF`���u���)^�y��!0[��O6���`;�-��v�<v�;�bǡ�`��3�Qvꄰ�cn̘���E����pht|FK�_�S��>2�=�g���1��l	�<~A
w2����(l�08��3`�U�">�OI�����kr1G�D3�(4��D���b�U���b*a��v�h��� ��TF�Eq�2*��PQ(4z3@7;u�M�y]p{{G���QT�Cvi�����H���ѯleV��r�?��UI�{�.���@�O�h�v��!���x"A�����8����|3�fu&]��{�p��������䗷�H�+,夑�����uD��l�f���t�c�䫦W{��E�� ���k��?�P��#�R濱�T�(�F!��wfK)��� .�25h������b
�92���My2Ǌ-[Ǣ ̝����>�6�_�Z�ϸ(��G��f�;c��Å�Ʀ$v �N�do�F,t�=iʈ3v>|�������3 �m��=ϟU��S�R�f��Lu����6�&�V5�!@�ͤ�
�dSԑ%��T�N���+X�=��`형�!�V]�&3�x T�j0�I9�����Eh
}f�a��&�1>b��C�ɇ��|�y������m�b�,��J�׎Y�t*I�U _C�|E�ࡉP��R����Z�[��O��Xطh�t�x|.j���\�db�d'�p<��%�F�飣'w��K�@A�IƇF&L�_sDj����W`6�I̹�O�%��.s���'anQ׃��C���d�w:Ƿ��O����������������
�!,+�#4�9�\32&JƮqr��jc����θ�U�*/��xJ&^�O�P�)�����Z7��9��Y	�][�}�fpT�9�8���I�!ċ+�6�!�!5���=qĩ����;�|���<�_B��R�C�=v+�r�:��$�;��t��5QX�+%����NK�B�YW�T���ھ{�x.��]�Ү3�v��:�eP��1�����M�����=�Ա8љHڹ>�zuiH�'u��5@<�e������������~�{*	{��ɚ��SGq+ʗ�RVpںk�t?
K��^���;�>܄<Е�媂�X���n�f�ťl�ƅ��Y��=�"9�o:��g�<��|(�O�[��A�L!����"7��#)��*���?T-Iq�:M��ж��������/+hc�a��:���>m�	uϚs]�����h�O>g��^Nu����.��g�!�T��=���c-G����g+0$Tg�ٌ6A�:Q��#�C>ym�O^f�ŏ��j6������������Ph9��ٳ�&�Ĭ��H1���u��L�ã��'��[��r7dۿ�� h�C���$�@1��a2/�l�����\�R�m]P��l[G,<��s/��>]7H���d���d4�G\c���p�q�|��k�q*׍�G�ԭ.�կ#Ɛ]�����;`���4�����{�#W��
t��n���2�Fџ9��ǿ+�?�Q�ؑ�:U2��|W�$�+9��I��RjA�ʳ�*�%�482i�e��x�)�V���4�ݗ���t�$/ ���_��&f�.�p�H��/l,leW�_|#P'Ox?����ꅏ�
_�m�;A������jq��V3jqcD.��W=��ֹL0`�����uQIf��ZU^c�^�Bp��YԶ��}�w�&%�������4����/�-��Pd�d��#�Z4��/�(�WG
�mH[���W�}`B�`]O%��ҏ����<�,z`��ob|v']/sZ�y��>x6�%��g��E����j`�%<9���_��̫>�U_�d [�QL��i���6�]��fu�$�dJ�=l�3ô͋��y��$��o����h�BW�+ ��N�� p�I�3���l�=�&A�;,q�#�`~loYok�>z���x���	�l�ݍ�|���f'<Aé�M^����_qߡ
�-h��@��޶O@]�Tt�K��������b�A�+�A�hU 1�MT2�9��K{��<ݛ�#P-�$:�}�*���ԺB��#=>așP�*D��Y����6��k���	�y�ъZ(X� Ӭ�����LޏV_,�f@���S�ͣn�ƣ���	u4���Q������F\����S3��atxYz��>�8)o���b�%���F첈]<�AOҷ�����OС�3q9<:1F5��`G�/�oXd����}�2qۼ:/��� �R!5� +� 1��ٔ�I�;VP��pǳ��0���퇯(Jk�4߷n�����lR@HC����G�.u*h5ejnJ"�NF~$�1ɋ�;Ӛ �4����Dr��;��&N�s;B&��b��WRpuѶ�Yː��'ji=�	�A/Šl�Y�r����۝3���=koe	n8F��G�C���J�NYk{�� �pi� �s��YĘw��]?���O�|m" �[��L\u�!_nG�=|ܝ�S���+�}F�f�C%����fUB�oxM_B�P�����I���s�Ϥ�n��9mP��k�=τ���_'}0�@��RA̤63&�$V�$Qn�����* �pk��pټ;C�Wr��p�O��.�
�2q?Z*@0Y���A��pI����%i�ᤤc�L��=����L�.WDS̹��
F�����7�U�[�lmXj�nE�9��Z����N�T�f$��-0�.u�S��3o^�Z��d�\�KY��./�~���{c��l�)D�׷��g:f�{4��?���EH��b&f	��E�3�G�^�2?͸w��w�����P�+v$�6�����1x47�+�X�lZ���5��$�ȰS!`RM�EꜵS2�ԯdf9�V}��_�]�����8/��XS�}Ѩ~H�fճ��<���y��)E[�w��\@S_>"xm��O̘㦈� ��~���i�Iz�2��t�1��PJ��6dPNl�Nv{���K����y�=���3��k������yucn�v	��#�.H��w�����>�%�뚭:��%��T��q)u�|�V��#����Z�������L�6S.,���jF�����.['4а��>��Xa�o�M��G��y�_~rI��\<H������ �<z�����E=>���S۠�t:K{Q'�j8D�V^s[Q�:ӫ�� �/j��d����F���hK�T����EL����gK��b����d���3	�Ұq�*�'�ٵ�O�P߯}?�8���#���
i�[�R@7g%�IQ�ϗ���7��%�����Dngd�	�9�QM�t�����r��:i�xEd�|,L�HS�"����;1���p�X���(��n��RD���i��/���$kb���|iL{��5����cL�'�T�x.��c(��ͯ�j���Gރ�΄��Tk���Xu0ǲLX�+�>�	{I��j׷�[�Ջ9#ީ;E�X�'�k�`Ü/w���`%�=��y��E�n�<���qlݐ��ʚ�ėq�.��6ݫ���`�>%1��y=w��ՠs�,w�0�WpyL��w�D�l�1z� 6��Qf���6��;�'޴ąj�Y1�*�5O�I�)*�o�n-������T[ �9ph�����\�2�/�=�SU&�@t���J|�Hq�y�ҧW�	���0���hl��F[���i䞅GJ;ߚ(�f;P��\Rq��uZ��Q��(	��ܼܕAnضϫP
�ohb��Ib�xI�W�ۓ����
�Ɗ_���F7\&��u��:�JS�5�6.dPc��/O⯃AȼC�B�3�C���ި�����\6'�xꃾ��
Ukq5�2�'��N�h�g)g���#��!L�[���w�J��,�~1K|�ZR%��(�{�R#%���X3G��V�ǫ\	�B��+}����'�'���}l �Ш1���bA�Fp��%'h~㉝sB�:�wcd�5�C�vr�of��]�j���%1�Z��kܫʐT����=b�RO��_ʥ�D�7��`+���0��`�����Vh���ǎ/�����k4���""�d���U�;�,�D�Bm�ld�����@j ��=mA�Si���R�����34��%�ŵ!�K�Г�ȕAa�o��>��y@�#H.�ׅ�6���q�v#���Y�9�E+��kc����U�q��`>$>g�
�?���6�ʫa�����]#�x�&�85�n�m2�\�8�Ѕ����F�vO<�	&-�r[��ՓL�P���bʕ�~R�_��32���tW�9r׼�
���xo�R?�3Hΐ���d�o��mH�pQk���g�g����UB���ė������q_"G���e�Y�F�8�_��<�7xrq�o�H⪵�F���S:����Ct|lG���h�׌a��rz�w�ؐ�6�(p��	FF��>���
BϢ�[S�x�ڜ���wG�]�_@� ~{�|qg}�!?K-��t�����,#�%C�D*J������s���h�s�K�g@��"�Y� ��x�X��,�F���N=ߐ$��D;�gk꜌��M*>K)�_�%��t2�~F��1�c��-b���z�t�n �@�9bP6�ɵ,X`��"T��8s_��ׅ��6f\te߰��:� �+���S17o"��%�hH��^O�J���.�OЧ7�H� j�W�	w�#��n����7�"����#�F�0�Z>����[��M�5H��.	��Jm��Aφz�|�(��aw�<oɴx9{����ZZ]�;������h�����[������D�*b�[�$����k�xԆ����'���˾/� g�7���a���)pe�� zz����f���Rӂ�;d��"%3�}�xH@��ַ(���[�� g?"�cB쒣�ӂ�5���EkS��ZAFq���$�T7��SL��G�AY�[�#�S��N�+u�}�������vwd�����/�C�*�����wx�U��D���yS�멧��7��J�/"�qR�u5�(���.@��&�s3�6�y(4}��Z����H�3�m3;��Ͻ_�X�k��
��L�W
�,l־�-̄����*�LRA&��(�)��B��J�{��}��z��� ���6KzS���D�3"�EZ�!vb��y�Maz��H���x]z@����U�Q�>�}��E��]^�� ?���w�d{�25�3�R6-�r�P�"��&44�M4?� o�9��'��1$��7��ٕn*�������%��p+���	��.'�SCEÄ�0	]�t�\�m�!'����r�?35�@�?�8U+=�6��G^z��Կv�p%�&���7j8~<J�e�&�Jd��ne���s�g�l�����t&]���V咈�Mх�綇Z�׶=+D�L(����e.݃�|�j_�K�Ϳ�BU��.p���[�(�4 ���N�!(���#F��m�E���]b����j����E�CT�ңO�|]�h�}Z��[�]X�// &�n�N�?���	�
7 �x5�|����5&뱰A��ȃc��I%��%�����8���\�T��ȇ��6��*]aSJ�y��E%O�f> ��|!��V?߇p\ʒ�@���Dr���B4�Vm�>G1��%�ܖ��

M������܇�:N[�Ofh��i��g�n��*�%�����ܿ�:@���.R��=��P,VSj����]p�m��;�1J>�־{��^~t��l<]O3UĠp�]�֝�h�|�02��V*��H�\�~k��
�:쟕�*[�5���8���^�1�<uU�묟�l��u1�kL���7G�����I)�]��{��m�;#��]o*.�X*N�]"��N΀68��ǀ��%.��Z�<�7�Ô�8
A:f����G�����D���r\�9�7;A9�o��;[k�Ai��ٹ���Z)�.�6�V�GV-��I�o��+?Sq�Eg���G�B�o����,!��� �~�?(r���C���&��RW_����i��u��l��ƕfrvv��pD����2�b���]���m#��O��D���i˩QQ+}� O��R�G���V Iktd�3�ito?ܤ]$�i�&7�,0(`�������낮p��q	�VY�j�=ހU`���ސ��A�oQ���)�*W?�P �i�G�>�M���4ms��-��,�1�0�^^Ɓ!����#�:~��8;�OozYZw�o1�0
�I4f��O:�]L$����U���P��^�;����װ;���%���e!��%��4��"l�g#���Ѹ��B��n��2�S�b��H���7�h���)�y�Ԗ������w����2��F4uĵ�ғ�4Â^��>�������2�����3���S�q�`��{��&9Qc&�}��v�Vp��_n�ۊ���?!�2)R������{��N�&��f@��0�c��BU(!��e��o��ՔW��x��L���z@Hb�A�C���HZ sy����貘*�vz1?�O���T�//%�eH���m��c�Q�A� �K����q�tX]@�I��N0�����ۢo���0��.{�*��xClv4������Z�c�Qs�Ͼ3�ᗐi�7�=�X�3ݘ���K�Z/p�K��.X\�+�-3|�-`���&