��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��N�]�?����U](O��q셝����>Z��f�0WK��{/���k(��i��]���5G�Q���_ Ҹ;�ja ��%����W���?f/
KI9���^C�r���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��
��?Y;���n�i�m�+R�����\�[���:1��2RE�D!�O���>í��ݛ�T٣��,l$��Z4c��XE�
*�a����>�:8�����}.�R?�Y�U�9�𧊈}�J��GT�uCn�8٠�1���ʸ�ל��m���"�JxH9�����������0�k�s��
\�E�LD�}m�lj�,$�؄�\�¨AYwT(t�ʋ�Ӯ+�J���/�fz+�4�c�`�,���t1���d�Z������4���7��I;iB�Ӽ��}ru�/J�L�:��+���%d'-�P.j�{"ά;�Զ>��,5���ýE^n�ϴ��&�2��q�޲a.�GZ4-�V�1J6����
��{���'?�[a0e��DY?6x3�ir��&?fT�����<;v=V��ƨɊ����y8;�R�e�jm��G�$C�Ź��K�H�=����#	:��J��U�FC���%w%�9�VY�`h;����3-Q`���dT� �!gg �"Q=/��P�U�c��%�f0���)�����I���揮P�y�MR�D�.�;�=��yM�9{����/oeԮ�u�l���z�g%�j-=�u��}C��B�N�W,7F�;��n�Si��M����na)z;q�u�(�$�W�+���?��P?�&R����Njր�(�\�5��>�ᶺ5�5?���3��%r`�e�Ee�tJ�惤|�H��IE��H���s���"çdZ?��ԋc��\����<�;����_�T�Ϸ]͊�ueM������=2Pa�%Rt���8�M �Q<�Z��kNA�� U�|��~In�;�&qpO<y���K�2�uȄ�����М�dD*�^CF�2��Oߚ�����ĩ��+v;�^�(��ku{�����SG��"�d6)d ,0���G�
6�/M��c�J7tX�/٬��Ԛ��`���+Y	�L�,csWCL{w�?s��zh�{��=a�9��l�f&��̇�G���3]��8Ef�N�!3�[��8Vl�~�zr#��\l�p?_!�F����yL�l�68�D8q:`I��R~{�(B���O�8ߜ����vbd�2/���aX������k��	�!�O<��n$$<L��f� j�-�ӵ���l-"�o˵�,4��~f�׶'���X��J����:�����A/�8I��O��#Xm�M}��X�)��#B���uN�D	E,o�y�Mm�ĸ�����t��B^�B0�[�1��d�[��K꼫���.Ȫ{������)��=���z��~"�5�O��%�I���+�B;�-�+�j"�P3S�%�L����l�ɾ ��݊�- ̦�?��/���$y3�l��U؍���6�n,A�T� �:
y�HXc�-�gev	�4�Hd� @�J����*Q��%se=�yf1�D�uP�O`���*�[)r~�X�x����p"�J�9E��'.T�I�aV��z+�Y͎\(��<)H8w}�4�(S5�۔p�0?�����ώV�7�BM
�Jӄ̧P��rKD��($'w��K�+"�wjhg�bY��G\�
�������K�n�I�o�9��\� ��Ѩ"+?�&�� ��K��'hﻥ�������l�ڧ���q���[�SYn��&�YL�8����Safg�IZ�0Ts����Xy���q0�u9�jT�~�)������O9�ȣ��o�I� z �<V���D�V�9̘)T
"�~�F���d����pi�֣�^��^b ?c��[�y��-��-b����騀�0+��~ְ�`��(ڗ�^���M�ў�q"�Q�4����e�a�*h�	�����eY��Ϛ��)�Dsz�j_��g!�;�����e���	P�`���#sp˻�f=ǒq�<8G�/p}g�/�'{#=]*P�\X�����c�T�H��̃�]���E��H�_��;���~�u�]��?��O��F�Oa���Z\\��~��(�5���{��� �pش׉���.
Q���q� u�o�mV�>��`�xͲ�D�g��6ǩ�L��
���$�C�4��-�/W�R��@�(��|F����2wN�7�#�D]5�漞Q���$�h�����V0�]ċ�qCK98�81Aҏ	�XOuK�U��d��#$O������ӝ��4Z�N��G����V�&c��66m�v��*�Q=5��K5���,G夰���1)�����W;@��Bv�>Z�Hj�G+(�"�"}9�&��٫�!(��婅v���qnCf����Y�a.%*4�@eN"�+b�.��u_�}� ]�t����"��|�#9�d^��A:��%���ϖ���"�C�A,�6X�5v܏�k�w#q>e��v�����.�H>��2!�V��Z�af}P���0!v91����O�`�$>�>��ﷷ��"Us�"Y^���k�Ɨ�f�J����ky��je�R���NOHX���@��V�0�� C��.�C���i8����p\��B��$�{��`�z�=���� (���1N&���! 	#�yUj磷�#�Wm����?��gm��Xo�!�핫�G��x}������k�\��n�]�kd���:l)K���{�@ڴ:��	���H�*v���s���S6|�Q�ރ��h��	s�����|h!Y��X��A'�CW�BJZ���ε{��wl�}�����4���Q	�,����/@:�)(��V]��-��^�q�>*֏��.���p��(��k��R�8e�1fUB܍�w$�_�Q��2;�Hi�/&W��5�H�(}��?8@#Vr8t[r����4Z������7F�`~���c�pٷ��|�B/D���+�pURh
���J
�uS�Hv�k�i^IkW���1��,K��E0��xc��� @O��Ʉo��0�g�B��m�S�� �I�$K剘��+Ư�@w'�t���
,$mW�ɀ�Ȩ�x������}]Y�!�X�~9.=�k�o�_̓ǆ`������෿�~��1@0,Nq�x�B���m8ǔ�O�D�j���7��f�Eo��]	���"1!2��~�t� nS-���l#)ݔ�qӨ۲3�߯L��������}1�ݎz��T^V�չ(C���V�t���29�����1/�����z:���]���[Q��'��#�J]U�WX=N|����^��L$�8�t��O�4"9iD) w|������z�S3��A��D��v�jL�h� 3=_��yg	�VE#�@���%!�^���4,	�@��f'�����Xozi,�"���I�	s��$;��{�{��x(�9�7c �l1�3e?��n���ԇ|���G�mis�q��i��[DLs��R/V`6"�K� ����Ր�B4�I�b8��~�)�p��O�� 29=�WP|H�%)��v�C����hR#��Y��)lGa��#	�����L=ԁ ���������p�~�7��#�(ҁ?��S�Z��k�*>����C��~���,F��(�QCx�'6�a�?�M8̆���Y�n����qH��^ ]�H<K����L~^��ڝธc*ux*
;���6�QN�=g.-��@O5&��ڐ#ػ%�v�K,�J�W�Da.-���P�yߘ��S��֖!�m4��i��5Rx�xZ������ڗ�π���$����k�m�sM�P�	�%w���B��9����5EÄ֒�K6IN�@�s|���""/jO��}����s��F�2�ل6�Ya�hޅ�~�n�N7�j#ⶦ��c�����e��b�P�50�fe���u����@��Q�OB��$�$�tR�>�i�-�D�&Fp9�(%��-I��U�b
s��Su/l(�"���d������P�U�S�X��_��F���(B]-q�,rpn��QL_v��X`a�1�hv2��ɭ��<�L��Â����e�h�ח���.1N걌l�z(+Ȅ��4���!Ѐ!&�o�T�TJ;+A�L���A}Ucz��]�
�����%y�J��ZL��C��vE:��+eϠK5u�1����'?q���)�R��ں81G���@w�7L:���+��r�	�3�c���#�?ܹ�ܶ���J�)	&:�ªw/��t����Po��ku���ɼ��።u)�@�?`r�4Yv�칰�Dxmvx텋�3h}>���A	���� 5���[C*zU�(��q�jE��@λ��z�b��e.�D4>a�O�?"w�|��#�E���K)j�O-⩗�t����IUW�����Se�K�7�l|w���b��V��g��)�&_� ��uf���ͬU�6^���z��{�&�J�)L���;��Gl��}��%]�uv���m�W��1/��+�k	F��^��t�-/S�2�N�w�Q��ţ�N��۾��_/~��ȒC~3Ӵ%��Wv�`�&0�LG�*K՝Pzt�Fu��/���T�+��*&�_||�|�B��aO�E��J%HK��6��c'*�0��(�=ؾBE��ҍu�Q���F|�CyW��'&Ň:Ys���m�U��;w(�K�->)5g&^N �����O�ƐJ�K������j��*e�������)J����W��V�C}�#�����'^m�������M�,��	��S��4��f��"զ�b�XdV��)|��4f�|���h,�]2�?��0���kR��Ͷ4�4Ut�l����`��׷gr^8��kx��L�`џ�R}O��)�WJ�| ����/A�[ݠ�{=����/����㳎�Xm�m-�~��PX��6�vy$��y�U~0#�p0��X-C;�{�2b@=ᭈ�uP5��s�
�[�wi33��fRh�`{`�)7O�5��P�y�ۀ+���C�VQy����7Ԭg}���������Q�<:�9����Yǔ��'Am���z0�؆��1�28D�,�D�
wI'	��<�ޕ~�6S�z�Գ�����f5��d�,���gwt�a�r����購!p���
�Z�WW�@6[wI9�LM��~H�ǅ`Tʄ��\�^.(����e��S����5���r���xw;3TXb1��n]�&<z��/?�-g����%Ē�L٬dq���>ཅ��}*�S�%�����q?*�~Fǹ�Z`��rV���65���2C;����}�R�?��!�D~E���Ǿ7����A=���P1W�R�̙T���#��������}���?:����r`��ٝp�;���^y_�j	��G<�����5'֘I��	��.c��o^��`D���
�OfI����چ�>X�'��p��H0�}KT_����Я^Z�#̶蚣��U�ԇ�^��*�iN@�~�<,��Eo�F�� WHO{s{�ݾ�-e��
��t/;h�)5���a{w���4im�2mT�X�ҞBA��5�6B�Y`��?A��=
�**�� Fk:����f&�4�6�d�ÉZo"�Q�+ lCogTֻȢ�Hf*����]���5� ��� X~k3�S�i�M�a�dB(ZB �%�S����wN���Z]�*�%)*�2�B�q#2Z��p �|~��ӣP{��,S]��ďᾉ�� �*1���;i�����<���`}��)$� �w�߂�'?R9o�����dN [#���8t�M�.4z�A7�H�jH�H�o�R=q��q'���Ѐ��}��|�<���n��MOμ�0(?�
������&N�J���v
�em���^Cv@�6d�
��Q�C9�G�����_6���*�=G�k�	7%��ǈ�-��ſU�!p#�T�3�`��m�?���g���� q>���x��>j,����xg"ŵFV����o(�]�5�g#&�H=���m4���Sw[9/���I��zC02:�bٰ@���in�K�tV�β���΅�o=M�dB�g�&���¬+\/Y%9��6�Q�OGe%����{�2s��[�������9:�}�_hK�n�xc+�zz�ͻ�J�����P��C���������4 �Im�t���7?v`\�����m�XbҎ�@��<��o@Oc�nG��r���a��0�<]�\�{�OMO7t�K�������	�`��`�s�3��bB���ܽ{�~�o���[�o1K�%�nR�+y�0#��*sNn�Ֆ�d]��!�O$]��ѕ�9���7���#�����Jv>졐$u� ��]Y�R�g�%���pØ���o/;���g��8�1%��_�~80[3˅؈�&�cd�W_q{�)o��^��u�n�B�1�(�7���ҙa�Ɂ�B���TiD�h_.Dt������{��j�p�1ϓ8v���g�L�㡘�Пa��څ�4�{z�]�E��[��h����<J�M�NCÅ�3����[Z���h���v����;�	��a��c�`)�윟�B�������-�#t�,��JE��%,���>)>�1�٢�t���ݘS(~fދ�-h��`�j�^!�9����,���u&�'m>XY$�Ք������!k,!S)��S�2�{��K��9"��"�߿��{�p��K��Kv������ZtO��'{���$(���5�y��E�c>)ٞ�j&��SA��d�(�(%�
^�`t���;x�ʃ����Q+ꂵ����5�-�S����ɺd�o<�Ga}��Q5���7�B����:
m���##��W���IMH	1m��y �s[�~o��*��p�J�h���u[�L`�+v}iG�p�l�x�\��Z�w�?�u�|U����MWU��4�9�7?P��ߩ6��мs
�jB=sa\����t��Z���#h�T��cFZ_7�}x�� {�w�L�W��������!@���w�r�3qa�8P�ؿ�Aޥ	��OBھI�8��9'TF�	F�>&�Y�@~�&`���'�0�������+�Аg5b��~�<�溜��=�JB&t�4L�f`q� 7��4{�qր��x黹�9ȣh�D�����=!���`�/X���寃 n(�gGs-�!�B_�e�D�P6%X�|@�![m"��XY��Ӱf]!����I���ǰ����_E����2�7���<%7��D�o��4�n8GK�;�5w 1�PT%��
9�$E?���5a���0�ڈe��Ь��V�,��[xt>&-������j�`;nL��Z�u6 _���/Ӫ��]@܀�9p.N \��!�o�'��̸߬(U�]d��Ɣ�CYf,NZ�o�yz#Љx�:��"ۑ�lT�Kͧ�Te�%�\=+�r���[eW�[��p�b#��k���6WzC�Ik	S��97�2�]ʆ%��x^�$��:'�ZҜz��F��@�m;x�����g�����-����n��ibc�|�
Cfk5<����!�;U�-�d�����4=��8���|3j�����e�Y�J��R�D���q���[�0X���5�ʵd��M���o�ju�������[��*R��*�s����Q$/{�V���hYuq���҅W���������)J��L�C�������N�j���M���?�AUPFT���Wn��'\���ی��b<C��5T���l�<@�ΨC�N�[o��V/��� �%U9�`Z�nJT���V��H��z"��K��53������QJ�����L��^��#��6Gw��
�Y@�;��Bc)�-3��)l�����H'�4' ������Pu�2�+LV@3����RF�^"$�X*)jv?Ȍ9+�h�s'Q�W�c�0���R]���`j��{y�I�I��a� �7�U������e�?వ�^6��|����b?hH�t$��o��0m �(�47�^����<v=�3����w��L��^�����7���<�;Vn=�c?�n]�C�bV�g$ju�㢍�e$=��a%��|+cP����Q�L�u;��_�y��zj�~桪�29�â ���V�_W���:��,1���B8%�V�<c�{�Fϔ���Ϩ�����qX�TN��o^�a���k=�^)`��SнB�����=�ϴ�;j]��w�@��%�p{t��p-�,�(N���*c-���4ϣ���U
l�U"�X��p�f�Dd�be�h��M���<�1fo�	sCҌNCX��}@T��芠�"�oß	�
��j

N�A�I�,��6��?ʘ;�9;x2���
��kM�}����(;��jMs����{�����D�\do���D �y}�/��	�ׯ+g�^���O��Q�N{pV��PF�ˉjJEߡ�H�;ո�(t�2�b�7G*pL>4M���M\�X�X��;xY���4^Fjڦ6��r���V=�Y���Z)�fTr�jl��I`*����o@J��Ts/)Da�z:܍�wp����
��*��Lj&�L4��ڭ�\+e勛qy8��5"/V��s�����KN�b _���%/�W/��ȏ\L3�$è�|��uH��_����;�y��2l'� �
����`;I��oC蟔������VƂIGQ�˱��h9��(ʗ��>�н���ǣ�R�������%�&���j8��T�XK��Bԙ����O�;$LY�
	�M���E������*�F�V1x`���[����%���Zۗ�����rB��nƌPY�V��lѩ���8��k��c�Pei:����� Q��^�bR�R1'��Ԉ��SV���"�����ss5��s�G�M�a��y�1pP��ͫ2)��A�g��8#�	�_��0��I13,�"b �z?IWB	h��L<�u���nO��j�*'h�h���Ԉ��gt�^U���d���><cjS�٦� �wr�k0��^E���^?F�1.��őJL�21B�^����-)�׊�@�9P��|����+\�W�+͌@���V+^�[	��7���gk��C4�̂�3S���=�ŧ��e��pj�/d=���
t	�{�<�%�0���0�{^���@<V���i_�p�-D'�����
eTH�C�Za���L���~�:��D����F�s�$�b�Cih�3\:�/y�L`��3�+�C�g�d��k�h��Lҕ�O��0bz>�Bط_���-ZH���j~��}(���;̼yӊ�)�+��̗��`�øӞ�:���n\���7�E�]��5��u.��s.�n�7$��;1ma�ܩA!��7Ѵ�Q�<�OC�1qO#o;݄�T��r����4�f������ �/��d�E4���j��6�P�w��#癕e�������e�`۬d�d!���2�E;/�}�a��:��V�*W������r)�B\�PB_4d D�����ȏ��t=�oaLV��rIa#E���3���n�J���>n=;�e(�F�1��$v�iڟ���+ֲ�һ��]��M't�T~��JL:�p�.��>�9n�S={-�H��3��ݣ��9H55��}�xjv9����ԩ�֗9��}7��-f���qy�$�R[ړĄ/�F$�q޼H��A�^!��kӭ���p Gţ�F�jBM�Z�5�����V���Ͳ8@�4h���TX�ﭹ������Ӭ�M�T���&�<=s��YI{Ӂ�u�����`�0ώXr,�JR�<&̧���b�ˋ���B�y�wˏG�_�F�v�������5���O�GtxW {�5m�-�� 9ٖ� (|�6W�����>�����,R_0w� ��HH�Ų��F��ߋ����ep�r�*�s�'��(3ם�t\��F��xq�������<��=d��sՕ��pQ�Υ ���jM+�:�-�E �L���҇����MMj���:�'��j��}��b�C5��8�(V,��S9*��.a�����٬�;3>WbY-w��p�DC8�R�������F9�����'W�"(#��X���`	:u%��ۙ���Ʊ�mD�t���/���e��C�C�HZlB���P���HY\��}��'����IGp<�#�l�"yX�'�Th�1b6�{�¸AA�n 3���ڇUj��-�:~Q6�;����J@&T��}:�ß.�y&�Ȣ��'E|�P�5-��ɕ���� ���i^�M&��+��7>g�$D�_"�	.�X?V�-�n�^�B׆�&���n� Ζ��y)1�OȘ2���[���	4
Y��@`��R.}qֿ������K+{���U���ɢD��
�$�>t�� S�����P$'-`Kz��%��l�os�A�N�DވmI����R&b�'�w_8�p�\�l�إ?�"����N�&ݿR����_�^g�����a�u>8W���K�A�[�>l���J��}W�F��w�8p��f��{�][#�mq���g
�Q�m?��e^er��z�d�<D㳄	%�$ �=6vjC�j]�>�v�8�>H;�"��H"t��$�=�K�=�U'��C|���W\OZܒd��Ƒ$�}�i�$̆�w*622��e%!ۓ�� �-��Y�3<ǡ)'l�<�c� �+����3��d	��/'@0C�sov�t^bMV��8��]���Tع��R���}ݗG|�z�1�6��لW ~.�>G�#H�X�p�-uY^���^�y��������o	}�f��N�=�sL8�:��$Őt�gTK���\��6��C�Ry�$Cq�*O�������C#mi�,?���Wr �(�kS܋c�k�� �2m��»��p�l��_���0�E"tK���5�&�,���>��0��T�C�'J�+e��L`y%	�2`o���BVsʀ�Q���ښ"�Y�'@8�{Sf΁�`	�cW����jmP�g���E�95i��_�!��Vn@���=!���x��F]�$y|�=b9ƫE�<�KI+ُ�H�Us�8��.����M;����y']J����֐<�#���"�	���y��j(��!op$��C�������Ƀ��.��v�`7���ڻ�� r�%¡���%�˅7k���8��pm�.��^	�^t�R،ѿ6rk��J��[2� �r
 �rg�8��Zl[s/�wZT�ϼ�I;d{�"��ޑ�����6򩨕�;���;��7�iN�V�"��i!#'S;�m7�{�<�*!~Ȭ���@�e��u� 8�����E]�ݑ��,��!��o�9���3����n	���T�����1��`B�i���	��jT��{y���L}����קr���i�j������4�X}��39�
c�8k�y@��^�V�lHT��I�!h�J��KR]P�=��~]nb��f�]L�m�x=��!^��D�]��y+�,�,i{�7�(Ѽ�[���k��{��ԏK,��B��d*�Kk�"o-�S�� �������ڭ;��GaR>:M�;IDf�����u��{Ao�6�������́퓨�u�"�R�l˹$!�mE�_k��,�Ծc��`��ᨲ1X��V�Il�D�ڑ�B�o�p���+�,#2��^��O�Yp�!�>��gt��N�����0���I��cI.3�dR�?�I���̇�V�U����-�ֵ�\�Dhݤo|ߩ�X��`{����dƩRdY�����n[j��0�����")禔�L�A�;�Q3+��� =e�ġ�� 6Pz++��;�r�U�G;��%ʞ6PS;:�n���EN&���͛�����hމk��e�*~H^�CR�	�=�e?/R��i.���;�P!�y-�|+��=rj���� ��m��LI<* n�Y�w�fU��ȱ�i��lн������tJ�Ko�+��?�z* �FyӐ:�@VZ�w���
�H�8��.%;����R�k�|)���ju�U^Ԝ��%�y=b9�A��)�X�����]�v� ��q�ja����m�J��+�Ov�B�룚�U��aߑ)�� ���o�؝�'<Z��,�'�>@ċ�Ŝ�D��%.=���jI�G<�	��,A�c�2$kWt�#��Óu��\=՜�h�������I�v���u����_���*}������nwH�IN��{���q�"�s�c�:hd�ȗ�v��kS�:N�zv�1�u%�����[i��F'9��\�����8(�Q�Q�GyCR!)�S[�]�}j��k5�_�eO�x7��5��p��s��b�M�t��f�gs�e�L�A��+b�N�};��`E�o�]wً;��\�3ƀ�{�aFT~��)��#u�����8!����*�l�5� �_���Sb��^����[�K�6l��F�x�[m�o�W�c�I���Ñ�s�9��@M,p�kym��@`Q��w'��:2J<���{���p������I.�s��H���d�k��������\G߯�8�SQͼ�KK%��v�o~�fto��Uŧk�]̐��"EKډAp�D�>����)D�Zn�����%��z��c̶�ք���33�Lc�|��ل�k�Q�����Ql~Ͷ���9N�l�
��R���
U��)h'MHtȏ��~$����W��@����+���Si|�>� X?���w��^ŶB)�:����,\wf�8/������A耘*��Evd�����$*�"t�� (�zܢ�OD܀�^�@�%��ƃ='�+��� �|0�^*Lk��6%���G�^�F���=, ;��S�B�{�֏�U��m�U������6�'s���o�hzaB��"��PSP�=�`�;Ҭ(U����}
m�}�ҘQQj��O{��wp�E��v�XT���@E�E��Q�k\��I��ƛ�0��7�%_x�j8:(���!�Qc�К�f�z�kaS�Y��gA��-��"���4���̪�ޛ��E���+X
_. ������W��"p��[��Ă��	�|�� W��x� ��z`F��'�|J�%�� �����3���;Xo�`��Ag�[�L�����x�� a�h����M8y���fGl^�}QLp���ɉ�4�D�H&��;���XS�:����7�Ҭ3�NL���K&h�p�*kA`����g -��y�:<4 �$��Y��A�+���Jq�^w��[$'�ρf�[1�T��:}S!�I��hLՍ���*R����K_o{2¼	��ڬ�D���ؙZ�y|��hP�h�/��,h[=q8�2�$#KZ̘R(l���G�gH�>�i�E_Нr^7c���D۟~
iJzh��?�Q��t�^Ҥ64�h&F�.ޞs��{��h=|�����Yk`2Ś�G4�ob�H"���)���3�<u�UV��u�]L�e���8�S�@�E'�I�-A�M7��u��+%��,���M:��l����zÚ;�N9����p��7l�B�NB�֔�n�aNW��Ra,-#_/�s�K%뚌��
\���C�ɞN郻������!FPu��X_VH[ M�����ma��Yca�}���E"w����X�>`�a�
��TGГ�rP��jU�uӲ��t����#ؔP�����5�7�,�AL���&�8��XS������a�e9��w:RW���(1���FͽFn�\jE�`�e�0\����,B`3�=	_�yNȐow+d繩�Fuo?l
�ғ�6�ʮ�r�FJ�sae ���K������qp�����?T�$aY��@�Ja2�*N�s�#��-0��O�J/%�V���k��,;i` .�H�[.;���z�93q-�z�b$"%-�qg	l3{���C�O�$s�*�Zmߗ�Xۄ|aLS8'[Pov0�J&�W��nV'�F�t�Z~��f�3	�qֳ�]��ׇ�.Y`[�'@}�Z{a�!+��}8�V��-�C��P2��r��#���o���G�ωy�;Gg,u�F!.�u?����h:���� G�1[���}42y#s��)�}�| �5�,��B���e�9י5Z$��T_�ѥ��>b��>ն�P�uZ��̍a�q�Crzc����C��G�fuZ���@�b��[��ϛ����\J�a��n�G@9�:%��m���?bq^�8B�K׽j�'O�m�Uœ�r$��E��l����O���������F��f]r��o
Ld;��,F��`?8�4�s���j�ul+߷�
[�x� ��B�y��~���:!ވ��&e�eK�B$#�DĠ��K���	��48�
�
�e}3P.$��S�U�kc��@�ؾ�OI����#&���H�,����x:=�?��Z��v1Jg������
6����῎��x%��Z�C��=��8��h�U�}��g�,}a]<���q���������,;*�'��A�q>��\`|�cg�E�3��X���W^�^�B��U���k�X!�h������j)z��n`�ߋ�#����8=��'��B��	K3�$*�������+��"H�~�h�K�-���}V���Fj��p�!S^B���![�:�p��M9zV�kA�mcQ��-�R�5�'�C,񲕖������W,D��*�u��W���&#Y�/�(�S���T$@��<��1��Lе�֪uX�q�C#q.��\����%1�Z�v@���"8�9�>øu��֐.K%β��S*�t��?�k���0�:ǔ�w��l��c��Ȏ]���	�]v��ں���a�S�,*��GzL�O����.�i�XQ�����j�$�|J�}i�.�y]��`rO]m��� �*8�l8�:<j�=�5?s�>�ݽ_@��y�H*�1Lc���`iX������oݝ��6�!��^�e�kJ�J�K���M6�]
KZ�nL�{�k��Z��*�|+f3�*AL]���+ƙc
�1/�P(�����>l"R�-�OTk����rDn+�\	E=w2�ӣ���#0��Z�	��JIP��(ٻ�r��fz���8��߫��*#��D����3�E*i�uwY]Iol��Γ�����o�־#t��}��l�9RW�ߑ���|�e@c���L����;���N��c�[���}�r�V����}�2����2I���hK0{V(�;%�G�G�.
,��܍2Y4n��@�P����	FԨS�N����� �W�2�o���-��3�,��$Թ�p�?��	X��R�$��;��K��$�p5���e�\��k$Y�hԭ�1�4,��|�>��M!*����
�5cT���$�"��5�V��/E�
'�j�� ���{�׶�2vb�l��X���̔J~*�l7��^c0�uS�I�⑆�����Օ���.BK�o#���\������:�3�e��pg
Qv����;m��h�77NzS�7�9HG>i{��#>VF&?p~�4������?���nvE��L�khg�������Z���q=��q��_�vn>��4���i���*����Bhz�ŧ�'6d�r����k���cqJ0�Ҵ���fd��X�rK��hU�q"��+�OR5k�ao'�S5Q=YE�|R�N�Dr�*(y��/Mŧ�^���3v4�a׺菑k�Z���R�����;�.� Q�G
�&��L��v�@��>��/}���TAv�YY����j�����sT��}���
����g݆��C�E`��bXRR��u�k���3XضY����c�!��z�{������x�㈖�\�y�v���q�}�隈<8�.�L�`���U�����8��u?b~�g��ʝ ����1�=oI���X����}+ݹ$S��k)�!��a���jD	~d���b��d�9���֗չ� �2g E.Q�EIWb��J19\�
��(XB����6V�d��dB
�V�*��r�3��dwle�����>�r$���G3',���>�c9 ��H�E/#2�Z�4�Li9��W3�/�%�Gc�6KePCA��Q��Z���9�Ӑ�� R�ub�rɖ=��y�Q��5'�N��[4�j�9��04����r�KP�V�A������Y�0ۇ��E1u;��uN ������USlf�aJ+M2�|�����{��o�U��;�NM���L1=�� �g����#%��{m�E��"�bI��p[i� ��`�9*��ҹ <�'%��LZ�~���${[n���� �-�Y%�����*Zz\���
'h�l3�t��/�d����ܠ��dk\��m�9fn�"!�D�D&ą�&��>��p ;�  ��@ �¡�[��6;���K����M8D���}���������7=�B��Y��*������ ����IS��9	�s&�����k�.<�, �"dt���EQ��$I�PI �u����FV�7�'ހ�3Ƅ)6p{�5&Yz�>',ix	�M����ۛ�zJ�r����-u�Ƭ`+B���	�i�&�t����|��V�j��RGO�?������_��$x�q�:��f�T3켧Akdr8���7=#������X@��&�M�=a�2��M�B���瀕�d���g{�Z����g�[�yFs�6�����2m�^-\���ydW��Qˍ�T��Y�M�i�k�3(S4mW.�"6nu��F���:/y�#��A������}�ז�.��]A����+3���W�/�Ρ㫹�(r��7s�TKe��"m�,�*{&qq"���
*��Т�0����m'g{p �U���*b�%�� >鲏�9E�d��������é.R]_CB)V�����T�p���J5�.��~Q�pʣs� ��=UEF��~��dT��rT��U��V8�v�������#:u!|_I��s�E`Y�b��=~���<0�5j�2Kn17eDt֍�k�6���W��.폇���-�������U;'�.�������8;P����fߞ��(ڌ0��l� ����)�N�yx�N���Q�i|N/%@��V�L5��|O!ivef{b�s�y`8�]��&;JOC���Q���6ģs\VRV�B�=ag���[N�ن|a(���U�@��Rss�����Ub #>x�^*r z	���[���@u�P۲���x2|Eb>�q�����a���rɜ^.��s@0�-��sM�`�\f��F�^�*������;��=V�\�� ��]f�=[7�qKi{��U�V$Z)&����4�
*����GL?*7j��W��]s��xI!�e5!�;��l�� ��t�v��Q��Kh!{Bd�r`��[Iȁ(wyn&4���Ëī�U��}�;��i�h����X'�m*�LY��x[/J�����=ePXI��Jօߵ�~���沓�X�Yy�5�����I&Ӏ:ak�i���Z�[R�6��s �2x��u��HO��v|��\BUN%Bqxv�X��o �ࢌ7-V�[ �sQ��^��!U���r�gɴ�n�q��ε���R��k�W�V���·������!��'4�,=y|w�p��f#C�ڴc�J�K�p�MmV��PP8m�x�a��CBa�=J��]� �/Qg�y�y�Vx�^�a��v>g��C���j� p��D��`�2*�SM� nl�yuSTWJ�0cJ/By�1yW�.?�F|XѾ�t�<�.�����͙:�C"��wsp}���#��a#������5b�,���)��@��z���ךv������u���
"m�8���Ġ[�����6Y����TR�iw���^1�M,�/���k��aW�"���9��BZ��2|��?J��x�R7�5x"�0p���u����'�GX^�ζ���8����j5޵�~7(�w)"bܛ�k�4�.�H�\	��(>1�Qt�в�/����g&����X�ӿ��(fQ���
��q�"-'#����e\q�@���P�ԕO~�3��fM�.���K`�{pv �RH�"n̔Y�ט������e@�y��%F�Ѐ4��Q�.e��i���=�d���FA�����)��~6Z $R�p՜UE�*4�L�"ɇ�Aڂj^S]��	�j���g'B��0<�w<X0RDJt�����`z�
7n���rܮ��d�r ��T5n���૙�)؄},�R�՛,-V�@���Y� ��w��<к��y�Cp�D|Z�JmB=�<+�ݳա��*-����!�n{W�(�\^��iC˗���ԡ�]%�������qF)a9�|i�<�nτN;^s�$>��~I��{ |�9����O3;W���g��ф0�u��;yo��5��=t���_Tdr�3�kr~�����:��ixؔ$�٤�E�� ��h�`P�!�o���7�E�&��N��b�ۈ7m3�E�U#�.���CҖ���TQG*J�B��k7 ;6�떫�BM�ܤ{���f'�A8�8���bk��R��I�[��C�'m�W��Uqr�HL���SV�1f�\5]f���օ⇾J	�`�@�>I_D��]?�͝���ɉ�eĀ�P��yJ�?uV�klU86���P\�NJ�Q>3�[���)�L�=�Al������=����|��m���z��|�;�JeSjpj��S�*�Z"A�*!�r�~k��~$)8�iMm�cKi�8�~A���ʿ��`�3�>��vhXtE����N�{\r�ObI���L6<Z,=ūI���0��4��qa�P�:&S��$�^v�+��x���yܘ0c�Μ!@	~"��� ��B�-����z��.��Ы�;���m�LA�i��&+ֹ4��	���֛�Nh8%ε���d�jo�2��ޔ�f���CTY�(���dZ�(�t�&�D��E���&�Z��6^�9��r~F�R[�g�/'�WX���(I
tĘJj��$*��z��Y��@&����f��:�j�wΜ0âM
� ���
4{5�".+�I�"��E�rg�`s8�]�9͇t�r%=�?s��4��`��I.y��s�J���!a�f���CIv�^W�^��u����qx��?�V�Q6]�1�����Lc��+�ʆ�W�
�����2w��^7�?��ǝ��I�s˼�W������ ������?���!��(�?սbWО�{�6A�+��t�8��V� ��A���ǋ��)l�4z
ݸod�o5n��*��-�j��<������e�VW�\�Gi� ����5R�L��G_9���	:"~{���I.S�pLO�6���^���\{��9VZM���J����Vf1T�CjS�i���9%������Oj���!f�dr�G�`j�"����8ړC9ou���M�ݲf;�g��lG�:�0R/J~	 EbN*Y
\����Ob
X
n��$K�>�\=�?��h
WW�-�B�+P?*,�
?N��[�Z�t������^��x�H�NNAh�zH'��zݯi ���1b�����.�h�+0�K����y7j9!�M���QB�q��>hp��'n�TH�=���h��Z�p{A"��0��
oy�T/gǷ����s7��E��
�9<��ޑʍ�Q�E2��Y_G;Z��}d(�o&�����[~z1;�\d~�N�9�S�{���_K��q���.�R��o�e�^f:�5���8�$�q5��\Ʀ���J�LOm'*�ˆ|(��#|�M4N+��G�V�";&�4L�/�7@�
b�e�#m���Q��(���qm�mTjb�a��B�m3�"M4���V��7��X��H��I�C��a|�փEܮ-û�Ξ&J����s�CK�MwD_�Ks��U,)_���ˬ�n�#zWj�B&� pI(5�m<o����B�h�^��A��նS����r�0���hUh$*s�H�����p���Sb����‼E���>�|��r�����Y4:�߉k��T||4��\�g�Э�c��I��(��sv�ъ�F��	��L�"�y�L�Ԥ���頺~����}N���8ڠ-i��X]�B���(�͕�$p�,��1�JB���@�����ħz�zUx��E�����@J�BL�:�߄� ڞR�e����Y��@�f*'��(ê����h�4��[)	^��hz
�Ϗ��Z�����D�����^nG?��� �*C+�u�qBY:P���qZ�4�>	�1k�M�Y�ͻ�1+��J��k�y��F���5p�V�9���_ph+�3��$X�>��0�L�ү}Ր�F��q� �η\�d&
���YO��0�W��4�����Y7
��:������-��\IS<J3�p�?���&�c<+ �7��}jM���[O�)p�f�򽃃��i�ߨ�<������o���fCK.97Uo��r��|J���������e8�>s��LM$q�m�h�D ���N5#���y)GM��RlK|���J4l�Ƙ�=>�k�^����/�P�[*|iz����!�:2{�K�����N���]z,9(�V����\�,l4��r�ׇ�C��ʻ�ZY�8��ޛ1����t�U���0��ΔfZ�
]y�v����Zm�Ҽjm�� `�}<��VXq�<��/Pu>�bU���%���{*�F����u�+���U���[�j<��8yEi�ø�A�,�����O.~�ð�͆ei��
��}� di���ҴLࡘ�%�(IʞPeրkb஥�9sR��*�;�J}p��f�}Rj髿4~�Z��863:���V�\�Ё�8�XX?�bbF�S�Ϣ>��9'�<���ݲ�����&gt��R��0�p�v̭�_�uYbo�H��l�m�2��b��[�ز!n�A�1H�|M� �u�6�}mavo��ծ;13���QH�j B��s�e�	83�7�����6O���aa�KA��q\n�8Na�R�Mh��!$:)a!� ,1ƏT[&��6]������z�p($rG��5�u�����
�M��u��M���E�Ҍ���Wd塎��Y���:\������(���^�:��X�! R�J{p�޲���h�o���B��tAV�>M�g1���Mi�1���{��&�-KQ
�6��ɰ�!§mx����^�_�����JO�E����7�������1���b�����6�A���ۂ��׭k7��C��~����u+�*�G�} (�	�S�9r���2��ms�
�3:�x��aC�^������k��b��#&�A���W�_�7���1}�E�e�'M�����D�a:�AP���M\R�/�_Xc�#�1�m��k]|�%��ݗ�Q�������n��i�4��X�<P��+IF^1�Fŉ���O�+9W����K{����T��&�`O@c�w�-��3o�pw \�(�I)0GA�?b8Sߨ �.h��-\�\~���焪�rCac�{�O�۠�{�t����m�Y�AV��c��E��W���$b�Sd���Z�F�K:�7V��Hʮ����̇\_�)��6��1��ݚ�!��J��4tH��3���\gQЪݳP	���M�c�1�\l�:��/>�6�L��heH�Z�7�}|צg��}�*���%	
]�&lRSz���mi"�'�:�3t��y�h���e���w�����:�U�j��V8��{�ӡ�o�R��{ն�lŬo���3^��,��3CE�V͍P�6YH� ��p���B�!C�r�`���Z�4��1�H�+Au���;��?�5��5�v�s���p���t	E�Y�U½���Э��#*���C�K�Ftp�]�oP;0�k2��"L�v+��*S_:!ސ_�0�"��o<�ԍjc�.�а;b�~m배�(T3�Z�0�h���!n$P�`�u�N��;kR�Q���W�iN��%��ޏ�{o��F�BH«��*06� C �b'�y<���W�HX�t2��غ{�t'��L9?�����/_n�nI�Ih��"X�N�֭�����o�]�*s�Zt���rΙ�ar��"|���R�S
�� ���|�A�ڲ��G�VY��lm
��T�j�R���L�T��w�0�E~�!ٺm	�س�N��o wX����"����U�r����w�5a�E+}�k�n���{���]�TZ��D_�a�`BH������=�H�$�>����[�1�I&�A�9��z�<���IK}.��DW�����	�}�Vh��4�D��0ѧ��j"��8�����+��_bؚ�EA��7�Y��+,o��$���ʧ��5sӋZ�㙐`RNDw�B�\%5Dm���3<|�C���#q����TY"���P����]�� �X?�~�¿ۚ�c�M �*��"���9�Z�ML�����}��f5m���Q�1'�f�-p�Npni��/T�%�:I�Z,JH]6�/�0�oY���Vl�2�|���Ў�ñ{9��{����T��j0�~����h"�FF�ܸ	A@��D��J�wA�9)I������P;��7��`4@z3)Y��o��88��>5ɰ��i�>�K�|�ѡ9%9��P�~�=�S�e����gf�y�ƒG�5U*-/�����g�sv7�AK�i���8�4��'�k�s8�}�����z&t��,=ǧ#F��c�����KӦ��If!��KW���^(�8N�a��D]RŲ����\�o�pFO��v\��DX}��঺n�sX�;�_��Z������n�X����#�/�:�d��F�-������^V�+y�sL+��3�BQ�S�\���c�~��k����ӆC;8=�d?��Z�"���@�QW�L%n�CdN�'�,Ǘ���Z�<Z���ݡ&��:���Ѓm���5�BR���c��C�:�k;��,�焽�~]�	\@J%5<k�3�&Mϴ,�c����,_ѕ�ٶ�bi@t����|�a���16��8�D��p���+�vX�[����5'{Q��m��n|��$����	�_,ȕJf���L*���c�N�q����^�ˈ/Bn��ѳgH�
2�
=F^d�R�U�{�2���Vҁ�+��;��Lf�b��M@�9l��eDԡg��M$�O��؆�W�+Y偑2�Wxk���{�	��9�@������r����pއ�+ܥ��F���fT�w_{^�J��5A=��S�.��;x�,C�� b(��@OF�oM>2#8Ul�i!O�l��Dp�N��0�}�����7�,'��!��8�Z���#�]��O�����1�8Hݶ�?�_d0̝�'��+�@YҲ_pʓ�n�Y�1ş�	���}eκ��|AN.�" �h���A��ǔ!pJ�!�Nff5�2w9�Q׊�$��܃�/�3ɀ�,zq��տ���b�8��n�-P��|�5M!���-��?�ٺJF)�w��\}�5�">��	������a�q�w�Aq-q��TG⫵2¥aߡ�x������"�!�f�>�SRY�H]�%I
˒���zuT�4ZGU=�m�M܉x��_]���0
���iC����זE���%�kc�k�l�0��۸xU#&�L
_!.�tk�*!E��[
T��+pr��Rnh��DF�x#d1���2�ѩ���j6��
��p ^�Lt����T��lO\� �X�l��xx��Xm��BT\=�0��f�'�fxAI˴N�#*E�����D��M �M��U�2���F���B��DŦvilz����֕9�:�M-�x,���g¨C�������ο�/��|ț��|B)��*������;mTb�?�"Lğ�����6&����<նΨS��h���\�_q���x���X�	���v������ ~�yuGG��g��,���G*�\�yn��5_m��Dm���fd1.�#2�%���c|)3-ڻ<����A5'F�vv�����z]�6�w4�U�)7���Z��VR#�T���w�e�j7.6����M ��)@|����~חMh\z[W�I/��p��S��(,���8��Rx�U�����!����5y����,7�
��2��:��us@e�/:D���1\5��8��cؑn5˹+x
 d�4�=`w5g�:o"�x����r��Me�Bd�O����)�FH��xzX����;7r��ǒh�X��}��u��|Z^�M#������Y�:G�J���D��F`��<q�V�."p�h8^�Ф�t�Ya4)ʾ\�"�{Z�D�@�����U�Z�9�77:�Ľ�b�O<ns�U����ɐ�uP�{�k�I��'���$HL̤����9����Q�_(7�M�3��jQ�t�#���^��i��V��T�Ȑf���f.19a3�⤰��6�u�n���,2Bc��U��y�́j�)|���<X��쏉a����-�4���s�9���RC��}�������HC��/8@�w��[d�v?'ﴷ/��2+' ��됋VyY��'��c��]7�àYƍ?]�1�{_�d�xq��2ś���P�؊�K5]�ހ]m��e�:�T�\��
͵�=!�'݄;���)cV��	��ܷ��SF�f���^·�fP����\0�@au'vxvg7.m�������҄�x����e�C�G�����I���Rzq��Z���j�n����ā^��ZI�t1�}꼀I7z���K��}�W��	?^���.�JF-����w��w��B��ZC��=���=-��My��#��n�ad�T������Vd�!bZCޕ���N�@C*l]�AO��E`��p����ϛ0���cK"z��>h�::.Mi��6���B���s�@���3�<����;�&��M�.�naQ�ְ_ٙ����z��t�/����(��BQC��D��n���r��G���
jW�E"IvtĹjW቟T��C�՟ô.˖�>�)-�n�������$F�\�h�"� %�A�g��1�F -��5ٱ�mPKzo�75�1�i|�B�iOp[�7�=�꠾�|���5���dʞ��F���V-Jqao5��7�"��%rs��	��3bk(�M?Z�ح]�A(+�P���BZK��ރ��©�ix )�o��r�Ui2��&$�,�M�w�����]Q�h���u432�������8�3g����7�l�-xq��d�-�;�S�3/���Dh ���b�*�V�����%e�}���]U�m�ٟ��A�r��L�`5�2a�qР�U0�p��/z{ut�QV���r�Lc����WD ���\>_���a:��^��|��&����G�t!{�o��}�ќ�$ğ���BL��m�F]�Z+�荢�\�� ��=k�C|y�C�I�,��Iz'l��#(�s�W9�*#��&��NҬV�#G����:f�����ִ"m��)�J7m�;Z�~!S���� j����A[��H��-	������@��J�R?vy�tI�t*4�	,iE�i�S����ѻ�N�*�rK(!�dt?8�(!����h`�"�h�\`�Ԩ��0����`;��j�,���[�L���L����(� \8�=�Շ	�1���&� 0	�RF/B6�Sl�MN"�l9�.�yɂ�=�Ñ74�`���K��^��&�"7�v��x��FLY�0\��(q���/��8������,E`>�C��� ���5kE��j�v���ڜsk���7-U�[�h�m'�g �ܚb8B���L�7�>_v�?���]"E��1�4��h�{|�~"�}0�9-<��B"���xI{g)n�\us�*U�EÚc�%=���$����V�X<���ٟ����p�>l��s�9vJ�%��V��!G�_1}O1�A�XKjl008�V���G �<;�㟢'�w�Ș��JE� [/D�ʁ"����?LJ�)��"��/���Y�3�n�c{cu^LlѨ@B�"���U���l�ε>D�O�D�����3�P/m��jeHv��;�����z�w�I�h�%1UzE�������"ȳ������>��7e+e5�k�L��#�<���h�3�k�x4CfKh�2� y���)E�u8���8��	�@G��S��fN��+/x��8����L#!���_�~ �a�@�G��P��\Q��)g[o��zV��(j�͍)	�-�tkW~��b��5jJy�1�V�L���6�x���~�͢3���{�6W��AůD�@u�6��� �<�� 9G/h�V�W3�]�;N�^~���a�I+{邳� �.��xe�����n|����-��.,M��dV(�	��%pɬ2�/��PN�9e����:���6س��KD�:P�Ӏ���L��֠��� �Ym��{����&�S06�m�4�%G���:��-�3e?�t���{���;]���%O��jY�Z�����XI�+�e��1��{��S�2 %V�{k���������a�w$���:���~�ع������>dѨS�[�Ë/��D�Nx�_x�g��n�w��;l���Np����O�@�)�S�ef�O��O��$Z!���?Qg'd;�ŇeI	��ˀfѕ[1����@&��v\��%pŋɗ�ʩ�hv>��@�̘���0���D/�v9V|��;L�r/CX�:�d<����#�D���FL��]C>ij#�o)��I��(�i� n��JH~TYl�[t��+:"�_��/���$����'�sM�k,s�&���ϱ���J�%�2R���fb�2�%5�֝åe�D�4�0�l��Ϭ�j�[��h(�������n�ġXX���J=e�j}bҍ���[[U�J����m��#�7���)�Z.¼z���C�|C/��gb6�үh(�֟�,$0��_H�Ƴ&ȈX�0$Gej]0����\��ߒ�w1�����X3�٨���S	ʏ1El�FvmFW �ݑU��{.���[e�(f.�s<��z���O���nO.�.��[B��"t��_0Z�%l�$zU5�s ���2B��lY&�؃�2�_V��"�צά�L�b��1T�-�d��?�!�t5��"�{. ���L6��Θ�T���oEHI5�G��uʹr��i�\�W��32[�����Z�k��pxVuVwa03^�.�P�J~9ގz��$����% ��,��#�`�B��Gn$*����CѧpC�
#%��7�B�ĸ��_��C*qAS�^B���ßVv%��EƔ�T~e,��b��<�R��4c��~���2�],I���Dư�L�
�Ilī�-���j�ܥW��Z��E)�E���k��'~�� u`%Z]�Ò�(Y!��w���}nlj+���h�f��������S��`
��* \��*nl���C-?1�/F���ǋ��C�i�h���yRt���]5���)p��^��M���B�Pw�w}�s�wj���:��B⶿O;�&�*f��ೆ���g�>��9����l���P��	YKZ�� ���W��"�u"m�)�شE��9h=L"t�i�#�ג�x8O�x�5�c�fr}�JB~;p �l�������p?osUL�-))��Y�vVғ��̞X~�M`^&u6�?�z ��b�$J^�O�
ll���L��}m�,�e:���?X�R��!6m%\C �1T!�p�T�Wj�Q�t��$^!
�f�L�~kcy����HW&F���^I�vɻ!C��?�w[�_<���S�RU��:&����i���5.��<y�����쥎�p�4E�m�uS���k�Z}1{�Ġ�аe�p�4��SS��w)>_m q�aϞt��ş���E���wT�X�5�c����Ф��W
�_J`��Z��OLC��L�h�^�4�rX��.s�gte�U�="uۂ��l��zr�ݺ?�mXB}3�^f�e�@U��a*������J�R�=֝&-�:��T�����\�F��?H!�Mj"�wO�;�_R ����B��JPDB�lD\Y0�a��\�m��=.�tst�#xV�Hki��zU�@B��>�nf�b�Q/2��3�L�E���]��D�iK0��=|#��^���ԭ�r%`�_~�~*u��x�|�-E,�X�]�~Dy��ujI�4Ê�pf,*�K���&ȟ�P��b�L�ݞ�+�b������01����l�{��m�,�M�����[[G�]D����0�A�p��J��hr�-2&Ѹ��,1� �Z7��|�fi����j�M;*y�� ��X�o���͑v}n��|��-��';^�?�M������*��j4��s��a��B�=�7p��X�F�뭹p�=���p�(P�H�g��u4+\A���+�O�,�hg`��&U?oc���Q��!>on�ߓ�-Bx�:[�-����GDc�2>����L��L6�ݺj������7D�e��fm��@b$�*��o�$Ġ��h`��7�G�u���l<S����BH����4�D=�Ζ�*a�^O�Ŋ�31�:�NBsh��`֓~��;��"n����&~���\�X����v��[�%�eA�Y���o,���-�b.�[�c�m�r+%X��3�N(B��A����m� 2^�M/K�8g³��]&1�h묓��9�1���qz�P��Ű�H,����R	�P6�'C�0[pJ<��*�e����2���`��
���'�������$R����Mz��A/�����0~3Zd^C�X���ݕ/#LY/rQ(���`5tط�WG�T�<8�+h��D��1!D߳�����%k2"!*�mج��]w� ���FqS�Eh_-�=U^s:��擰L$�>0��ͮ��er?Р�sOR>.{&޲�o����l>�@��Gj��;ux�.;\C��� �Y3�4�b2��J�a����\�<L	Y�����$ni~8�)y�<f��5��&�Xr����
�I����U��g������vr��g��J	D��xCh��w?Z����0#ɉ�Ä59j��A����!�A���⁋��5�+Ղ*�{��wA�Ȼ-�S�n��A�xF.r/��ưG����M�:4�w'o��l�/�B�չZS~,s�GϤ8��GP��h�?���-y�i�}�q�
I?�j	Gu�*�B�?��_�+d�h8����vPH�����q��mυ�u���L��l��R�18ތ���F�ᐸ�3�AK�~!z��'�i��4�54��A"��P�՗n��2��{E
 %���hT$|6�6K�|)q����D
��N�y)C��4��_W�/` �h,n�u)�-�*��tK$.ہ�ѵA��Ï��������R(�����AwS0�u��p3:���|�x�퍿���=���T����ֽ�cٵ9��3��>:u��B�P8ړQ�s?���܂���w�CGS��isp��`���x�P�,�O����t.'~��@��+�Ӝ�c40�_�X4MmU���\�c:�+O��C�n��}�`\@_+]��'DJ���G�7ʨ�4�r%ˇ�;�]��[�i@�������T�f���ʣ���A�A�U�s\�/}�Bz�sk��EK����h�s�Y*ׯ���eq�Un�_��V{�[ђ���� c�r�i�q�C}��/A�H�k��<�:�͏�^��d�>����~�W���n�Dt��>Wg���?Y���<�Lf[JR�؈A!��/��� l. �б"����u}�(���v�G:ui����X1���G���G���n�Qq�� ֭�@I�H����&��}U_�B�QH\'`a��F�5�|Ý<� 3�=�u�N
2g�����a���D
2r�}u�M���M����ޯ�n�T��n���!H}�``�y�T���q�}��ײG��g�p��r��cxW#���x�[Dzc���9$���t��%U9������.=K�H�Ka�����GQb �2=4z-���l��7ZE��RCc�@�B�CB͘k�D�l0�(�Mm�2�pI*����ǚ���J��셡n��a�(k4�f4�X�ן:�Ҝ٫kj��<�ν�2-�7ҫa���x��g�D�V S[7U�OëVcȐ⼹�����T@�'iy1���Ø韒{ti�~�mi&��;��7�U.�N ��=UU}�9��G�������}�K�to�Ky���:I'+����f�7!%ORe���������O����N�]:*c��i_&W�PJ��?���s@8�!��?����0�_��������Tp SDl���MpKJ�������b7r����Y��1���J!��偭k�o��5"� Y��gu��A�����$��߆}/�J ��$�7Xo�Z�F
����B�U�)l�U���	���Z�5'���`;4JY����B	�<�i�����}�˵��:Y��nNȱs!����0�Ok���K�O��0t�z�,@7���_T�`o�K�K���N� �X�rsfy���iK8��3P�΄�R���0�ڳ)��c [�W�G�<�/!��K�X��\-�K	a�YZ���4RQ�U��nl�d��6�OlZ��U��t�����\��
���	��k�j�L2�f����(��iN�w_����h�Y���b�����IF�J|�ZJ��y��i�r��( ��W�8pL�_��|�՚����\�sL",�P���٠�q�Ώ�� fIR��j�[�ĥXE}�� ��WGZC`�$Lխ��x��'�|��]�.�u��h�^��/�<(FF�B��Y:��p��L.�?qݑ��v�G���,${v��n�;^������s��vh�7"�c��Aǣi�H|��\�&��6��a����{}Ɯ��)�:�}#������H[�_@.��53�K����e �WS��=e�S�۷��D�dH<+�>�1�I�:���;-��X9y�٨cJ�`�YZ!�4H*�֠@�K�3Jh*��!ƅH���W�O���u�����@`{�k��7wE^����]j�t����aĤ� �a�^�B�% x���O���c�r�6��p�R��M�7qMc���h��,��{�~$�v���M��:�L5'�N��iV�������l<,��E�M�Rrn����f��dN[��E��&rf�OL1�G�4(�M^(��X#�y�5�����cWy�M�!���#�rI�7E>ZGRj?><2��q�ٛW�7����"����N����t�i���<��6�����տ�و~y��������,��h�&s�Q0���rP���`@%�{'�F���GQ�����8}��-5Z����g���N�|IK����?!f�J�����I�.�+$Z������.��[��'[�"hK?i�蕊��Z������s:vT�腪j�\��5D���?0k��X�XB�%��C�b�ڷ��B���	�;ph��r\O�<�4d4:�����%�9\4~��?��LiT_�	v�a&7"�n�vR��pXgvI�W�X�	IP_:����F�%��lۗ	�5��G��'l�`�,�ɷ�R��P�Y��-�5Մ�䷓X�i�a�+��6�x�_��Z��{��u��!	K������L?,�9S5���H$f�:M�k����&�żJ�B������v�C�.%��$�{�E[��]�8�Ni���o�70,gIa��wSE)�Z
�ezK�|M�k���@尒ڰ��D� �c4'0*�>�ݪ?T2Y�V�����s(�z��� i�#;���O���n�o~�e��[�"����U{�!j����Ù�Opd�F���[�rcȅ;������-jxi�AQ��*>2Ӗ���a�pPg��ab��a�4����!B�(�|�ܵ�`b��'(��!����ȀT�9�)\�qΆ�'� ��2��f
��s9i������=��8�7�@*$�~!�T��K!h�bwSژ�ݣ����P˴���F�:GA'y}r�ti&��z�<T�O_<|mz�M�t9LApQ�ں�C���?�.rcPN,Qz�m�PV�=��o$��d��Y�����
�����7����$���KK�8[tڱA�*f�a �[\ߠ@{z��5+;c��*���
K\[���Z1�L�3
POR�C�e������(Moǟ��Z��t�ٍה.L��5���f��g��_4{��^�&���9��=}$�<����I�Q��ΰ��'�/L���U�,\�����N��n�������-'Q�a����U�bC�W�`r�(�q~�![�?
�0��l.++�5JȐ��8���x��aG/��Πc���N��I���֭�C^/ZD6ԫ0�
�
X<���J�p9}P��d�>��aؗ��.�O�;y�ЊT�`��L��,�"�r��I�h�L���#��wƋ��h �˦����� ��s��'�@�~���Z��X�q�I��Ԍ�L���X�`���*�4��Z��S�#���F���!	��:�T0�x��n�mQ���v�%�O��ߥ�'?\n���t�&oa���?n�E%c�)�yڝ����*|`z"`P�Grt8I:>�0�Mq͙�bt5mb/^��=M`�fPW��
5u{-��$��3��\�D��]���u T�&/�Y�I?�G .V�glֽ���H������6ϗ��4�'�PTiͮ6Ë��5�=(����hx� �ݳ�6.�qTؓ�B ?��p������Z�m?8t�owך1�ˁ���Vg��Yu�#�|��<͏����0=�ѐ�������pƎ�u����@h��
���Ü��%.�/��*޺b�Ͼ4����g^y��<�Z�y�[p!�&^G��Y"�/���
D��@��]_ے'	�2o
�m���EBK=D5���B�Z\t"0ޚ��m���.~�� n�� �;P�&��)�IPa��y��1-�ܵ��Ux��1kJe��KϯԎ?>���	`���1D�.�m�"�M
��n�P���A\�9M�⺱���d�~�/�z��e�7	�
�����������HK�a�Q?1��i��f�(���"�Z�_�\�CN��K��G�](G� ~�.��'�+�B��I�@���2&�G�����4c-�����I-�"��6�K��q�~��f��uuٙ!4�S'�s3@�`��@��$q8��A��xn�9Ӂ�$�6�b#�CGJ�ƙ��_O��V5�O���?����.�r#��Ţ�1%� ͪ*�Q�R���5�b'n��1����b���R�C�Q5�m����^q�x،V�Y�ﻪ'�����6�Jd핯<S�����7�8����]��88=��.%?V� "�RK�.fN�9L��T�0��%B��:t�D0zMD�0A�-�R�O�Jr7�{���o��,5,�.�[S���j�4�h������1�W`Eѿ��4e#^���H�K�>Vk��3�^z�yK������gy:7S�O�3Y4n��l�3�x�q�����Ҍ
%�.��>�Q�p�e��R:R3��sq�- ZK�M����z�=.-Ҕ�/��2u��<v���ϱ�O���A7
�i��vA(JE�U��>9��cw�]`ل���������oK.�q�V掛K�#\�%��%7J��s(�A�;�c� ��M�g6��c>�F��O/#����v�7W�����-�'+%���z��E��_m{a��4��z����x�{��	��.��|���.���O�k��-���8I���T�4x�su0�Μ R��Q}zfeӝ|�A�M����6-�R�&x�����
z�m���fG�����9`f�e֚l>T��c���n��#~D��o�%�?)H	���PFs�;|���7�����D�wѡ���m�o��h��P��lc�4dd��I�0���y�2�(����r���b��Q���p=��>���жj�>���!��ږ���x�n�5
j2��
t�9=����H���5��?�w�X!��d��?�#�EV��sX���4��Xt��^c�&��e'�/��]mm"d�B�Q�\�B�|r��a؎��+pn�-��թUq�W>#1+�E��8��@�4�5Ǻ�N� �vY�)�����eV(�r\�-��a`���R��/qEj��)�٭bOT�h�XN�:��2��ӧ�J�mA-�/�l���U�e,��Y@{Zl!�c���ċ?!�:�ۣUD�O�cl�%��wKO!��˨�藄t7#�'�]���i/�~��ZΚr�`�i{����w�6��B�	��������J�Kv�j2+:J5�:D*��!��E�����+�6EC�5���u�j��A����q<���� 3���I*� �=o�߇�\f����G�_��m�҃��el�My0�� ٯ�T[8м��,Y�M��XK)�YY�F� e�hp��QXjR�d(���W��Ha�
2yO�~Ѓ����Cڽn-���ղ�xv,t�Z6��Q��>�kj�����Kf���=t҉���b_���I�wL��w��]����=��<O=U��x`�m0��ĳ�#�05�г�����A��d
�e���H���
uqp����6�@���3�j��]&���a$gl�S��Gj�'G4״���.�
�'�m����w�k�;���t���S�LF9��רbH�����W�����N$����*R�[���jq?Xj�W����Y�
!�tSz�P�έ,�=�Tǎ7�m�zq��c�X?m���>66�G��{.ڎ���b�`�|�M��zQ0��W\��)���&j�����p?!O_��a�{�v����'�?��2�p�w2��A3d���c>X��r)��7V�1D(�w#E��Z&n��� ��u���ҔQ�z�ug5�p��'w}V6jL��	��*i�CZX��+��S�'��q�$i_�e{��+m���|��K�A�ƌ�LK؉�2�h��\��`fߡN��3n]��&�@���E�����T;k�����A:b���b�_�RU���qg{�4�Tw�K���pĩ�mI�X��	s�Z�����$f��Ã~�59�/��ugo�nA/H��J"�,""l����YNBm⪃b4���*x {8R2�#�LS�
�귡�`>B4조Cc�wf�)H ��,�x[ի�W�Ku����m}����hw8!1�z�"&��=�6�vW��=�7@�4�0F�����#]u�l��.�65��}P,�ȍ���yi[�Ŵ�_��td�s�F�o0��pY�<[�F�.�\S�&�up�8�fa��9Ƃ=0#�m����� o�T��h��qY�;�d�uEXִ��!@�p9(�huuJgm�U��]]���;V*?��W�+ ����R���twx��Uy������6*d#�ӧ�i��^:�q�]�m˛S��K�r��s��j��.� ����|f�)~P�r�Noƈ�����N�;��}�RPps:h?lM��?:Y��d��$��΋���s��&.ɲݭ���!������X'v�$̐�B��Qw����_��E? ��g,��
�W�����Ocf��B�V�>�Ixٕ��&�Q/�A�c��\�S�'03�C�9���~bH�"��2�
Uo����-������^��LxR�����ε��R�
u�ޡ_w3�9�=O-2�i���E@��-hi�:k�⩚k�Q�?Ug�,��ga��g�;`
�R�MLwt��G2�9�ID9$\����!�M��
-T�����ЊC��Ax����}�]��f�H����~�zǴ"�m�L�.����n��&{<ko(0I�5m�G���_�M�M�U�m3p��ʌ�O�"!N@��RqؼI�����p[o���؂o��5�s1��U�2Y�3����R�8:��߿�|��%��3�Xl �,_@+"o)���i�+��]��߄e Ɍ>ߋ�w�^d�M�r����V���I���d���q���m;4CK��7��:m���i�ޭ�Ν�#r� U��i�6�Ǥ�G�\f����z�O���1&�
$����z�N�l�Z�|�k�W.!�.�TR� ��*	p`5((����Z[^�Ub�M�������a�*��_��3��Wôt�^����k�F���o1�{�E(U�5�$������[���k�Q��N�)n,���2���M�.E��cXLi�wSka��ȸ� �O.cp)޸�Վ��Eؖ@F�����Nѡ/�#�uyzE��K$Z �D��򅫲쯄���N²އ6��v���G:��_Z���ȟ%d���l�!�X�Ч.�����j�C�n����1��"�w�JF�
�ǩ�����0�ʵݻ]�1�U_;�2xV4�v��R^.TS�d�CϧY)x��ߥ±c�YJ�2q��
#�t�
S�7^��'��i�f���{�i��|ޮ�	�G��.R�D����v�l���Y���ud�������Թ@m6'$���uz�ھ�Q�ѡ����ʿIO�3h��(0Bi����>�H3,�+f��m } ��l����gG��	�$:LL�]0p��1=��CG %�W��@A�lc�p���|�]�]Mn�x���@��m�a.g�`��rA�qw��]S�n�[�%��ρ�W�N ����KwݮLK1^b8�?����(ag�B�G������B��k��X>�a���RG���O�ܡ�2�q���u��(�mo��<wE0@�hlSx���FzfZR�>I҂|(��*���ǴR�V�>��ވ���[���U��֥��G�p/e�8Ϥ��L�ע2��L5��c���v�i��<4��̶bk&FҖN���Q��N�������y��:\8*1�9>.��1N,$��<WC���e���*�_`���D��u�#�>��Z��� �$��|����['V5�Tu�N�/��)��ט��Mh�Ǘ�Ζx��p�h�f���1� 
�שļQs��Ϛ�y��W �_B^����aN�1��ϱ�9@dy�X�]��yy,8�l��~x��qQ� �k1�6Hw�{1���<Gm�<���F, �\7�ϰ�e�W����&2w�������85�{��_�\6U�s�,F'��V(g2������3#�?ȉ�w<���v�.�4�k'�ۭ=S���'����+om,�?����*l>�7
������ɷ�� ����$y�nJ��yn�G�R�,$�K�X�\���{��z��p�@F��D��Q/�����nh������@S�d�!�!���Ć�{$��� %C�`��N�Kk��,���䵥?*k�h�<vהm:�m�֥u� 8�c��B�*[��"pC�J�o�k�}�h߸vL2I%���������$�7_G��d�����哵����)D�D�Co�~��O��n� �x"�1��Y@��b����m@F ga�Ѣ�k�h�a1��og��:_�2>P3x��H)xO�ڟ�kh̷0R>���*_�A�1T�ʬ�/ݤ���*j��~��Ћ��@��������Am-�V�֎�(��x�"�:���J�횽�ף�/����4՗���Vs��vo���5:�,��A�"~M��SR���Ŀ;
*�"�pY�2��h��KxDd�y�#,�B~�sܔ7V�ք��K�~�U!dGQ��SAf���c����+KZ���D㐨S8Jp��-w��glV��%�5W��ú��!��Ӄ��L>�0�+����z��?s��f�!� 9�����yr�]�aɈ����q�bX��r6��W��׏[R��'}@�O�m�O�@o�p+�� �D��re���i+�eӱ�rYad� �μ����]!/���!�S��n�]ZR�[!��{������=L<��(���g�<]��i�g���jA2`��V�.�Tn���=�Io��cij����ȗ"��o��Hc� 0���3�9��[�19W�6.[U��]�u����Z:H�H6��o��Mt�27��D.�J�cI���apkر��$T�>�"��7w��)�D�Z�r���ȡ!��0$���e5�$r�㐣B60�8_ܦ��i�Ny#83�	OX�3���
������";����i9��z传',7L�/��HK�)���F���#7�@��{\�~?(��ݔ�	s����@2~�W���5�X�q�I�r���"@�4z��mܞ ����e,gȀa J�y="^��<��,���.����p�Ɲ+\4��{5ug`�*h!�lX4������⛲
 _%D��BJa���S���f�+�r3�L�(��|��f8����?���[�{��I�XɳBK8�$���n�'�|����IA�
$GE��2��z=';>%��@x��!��c� ��{�쫕�n�\s��"&mm,Q ��7隝�S!ȿxƟ�^	�oW���"�XF��FL-�?X{"�|��)PL�]�*}��~��<(h�25,H�J˰N�t���z�sl����zD��I��w»f��&�lK�g	��[vX����FuF�Rꈤ7�{�ak�%�s��(�wc�(L�T���+9�1�	aa�E鞵*b�`�$�~t"K�=F��]���<����U{�$Z��$Y��u&�j:wלA<��E��Tg �g����5�P�k��\ޫ�y���F"�8��Гm�?S�L���BK�4P����{����9u׍��ã�!A6��j7�9���'����C�|��]�-kZ�d �I{ V�%�D���7�����G����.W?�$˃<����-+��J��{�)����<Q�{���kk�޲�v���yV�_0"B0�-�"��0�YR}�>�\��[���ZI�6Hj�Җfv����KE?�IR��G�4Ш�0�Ծ�:�������������5
�Ǌr�� �o6�Ÿ(+��$jپ=�
�;&�̳���f�&�vɾ�>�42�^����\�����p�.!�(t�W��.��/�xj�)�3�yU>�����0�&��bj>鐥/]x<fW���S�Ϳ���~��W׍e>���I6\��������jx��HG46�����<*���wH�!�%�7ܱ�H�7�CYζ���:��{c��(��`+�~�U��e���R����i��UH�����gQܸ�pڕ�]Im�C���7jK�"kPL}`S���������`Bn�/�jo{:�~6�Ī�+�;���W�~��u�^9��H:�Af�w�g�UX`/���&+���s	��NՇ�)�t�O��,#TmY'7�:$j��r�ǆ�}>�����Eg������4%k���x�[d��t����� ��ìQ}ߝ>��Vlo�VY>��0VB%�I�\ѫhۚ��}5�_�*�x:�Ʌ"�<��Ly����[â \�������ZщZ���0�Sx+.�hO�m���7'�
1~L��1�~�Q0��K%��Z;��IZ��S܋]�[&֬�h�5�~�xF�� ��=����TخI�fYtG�A���_s�N����R��T�m�7Ж�Nr;	�f��	�b��@���=�7��J��o���2 X�Q��8����4V_��$2�@y�� ;Ȉ��TTނn�������z�*�	���O��z|p$&��L|��ղ��\$�V����ӶI�Qd�rn%�Kj�0�d�2%Z_z^�Ӫ�-<x�;�I����H�=6ZkA�5?Uu=�,5��������Ø� �^_(��9�R� ��d��Nw��z�2�#P��[e�i���d��^+��>fI�.$+�xR�,7�2�4|J䌕�a�rҹ3��dL��I���H�'���8A��8w*���_je}t�m�����6` g?�>K;o��.ˀp�d��-S�� �P���Bh���:��M�?��i�����Ő}����*���VTl���>�JZ� ��aߚ��(��5�H`��� l���=�ޑʽ�H�Z� ��� ��l���f�⊷Z^��4$ V,�1Ϣ�4mXdI�0��u��
����=�QbR\�5 81��������F�d�a�kp�>F�66��B/xl�7��Ր.,��R�v�Wdw� 3��4�;�<H��tT?_D�QZ��T\�pW ����a�Kw�p7�kQ�_t��W�-6��tg,Ń����.}��4	�ޕx��G���(,�u����.�~"oy�^�+ Hl�B�\�Ȇ\H�B	ƥ�J���9�M�%;�i�} �h�y�1��2��ץ��F��[k�t耣�@�6��,�%c�����* Ng���r7��1L"�d��5��%�s,�	p⒩!9�ÎQ�//'�A�nw8�Q��3��:�K�K ��e��D������@��u�L���Xɛ� �'�	�/`��t삡4br�O�xd�I��m�*k���b�ٲA��Ѳ������ ��wZ9��$2N�x��t��9����a�U'f+N��]�}oxpbH$�a8HC�}�³v��MWa4��ɎY�2��y>��Y'I8b�!��q�R�4jqpHK!����!LFQ�͵�o�fO��i�4�/�)�P�f2m���r��~ph�Z��vVe@�[.7)��8������&cfbP<R�]a��j�ŀ:�����K��XH���0C�1�B&�VrEwj-��lƀ��>�3��]t���	uL~��`��@�˦H@v� FX�q`����������y<�1���ٸ�km�]�6ަNBq��`�1H��ȅ��af[8Q��+�I��}�b��Cq#o�D����aȉ]>��9V��H�d�mY��ڥf;�f��~}������ /v6�=��.�tQ��=����q�O[�)��΋�`ͣI�;���]��F � ���@��F���5�Cp�<��h������Lq� ���/�r��$�'�oEF$�}A[�+T���*挃�� \L7�������b's VIk�r�f����J��v@Ϳ�߹���X�2��7��=Y�/��ۑ��Z:�[7^����5O4�������6�ͻccDvh�6�E�N��%�}d�XzLl0�0�XA�!�)h?�� k��P'�w��
���Y)��V����O� qr����j=1ޕ̴�*���t�/�|6ޥ���:��e��+M��v�S�lknv����l1\o���;�z=��ϧ �H�_Ѱ$�D��WT�������t����,�|�qmg�%��-��
��8�C�,I�'ns�t_�FR����(<�"|�������z���6��p(�Z�ԄD�}�U�b�b����*��L_W�?�3k�C��<��ۼ�k���O���L���'3jA3Y������vγD��Tێ��� � �N�[+�	i�Ǔ���7�_[�@����u���Ғ�LFFޜl�C�v�E� �ǠfV���S��� Z�y���ʄK� 9��A*}U�I�S�����o��C�4�-m���m��xw�nxU��˰��E������6���������c(e�@[��"�Y����b�ۻ5�� o�,ƙ�I��g[�M���Y�&���T��Ò��=�p����T21�߳���P#S�˞�-��a�4i��m$��$�G��ؕ�aO����kDM}	W˖�{��'�,����`��w����Thg��|����;8�7�(���C�KBʟz����ՙU�w~`�wc����{5�=� �a�U)�C����N��X��ެ���.X	�L��]��뇖�m���_�M������$��v�9��.}�=~ �`7���X#�Nأ6p;�v���Ϝ�1�H�;��P�1q:A�H��Y��%+���F�r�����8��.kq���D��2rׇ���Q�*e��i	-U.ʘ��S�|�P�86	Sp�w��I&)aH+>�G�f��5���|�'{s��(���b�������z>��b��\ݧ��T�%s��1�_n-�B