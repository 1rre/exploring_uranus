��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��N�]�?����U](O��q셝����>Z��f�0WK��{/���k(��i��]���5G�Q���_ Ҹ;�ja ��%����W���?f/
KI9���^C�r���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��
��?Y;���n�i���И�A"�vh�?�}_{������=ٕ;P2]�k��ޚ:���,*��e������7�`�ק�*2�`��ǌ�Om_Lf�Ͷ�;��AI'���4@������^�
�:��r%��<���U�olt�9��̼�_��r�V�����y�������N�L:��X֜�~x�<,2I�`A�<
��O���� �ȋ�P��7���W�iݗ��)|Q!<��ݖ���2��J�6����������a��g��_���pUk�R%Ck�2|��mJ:���T��BR�k�2G��Ӌ �(���]�8z��[���[l�O��@� ��I�\lV%��j��Ԭ�m���s�TY�R'.�%Kj�Ng��a����������1X�'[����>xѻD�'��J鳩pBӭjͷM`�����ѰE���C�[쵯��{,��q�`�Ye�!�7/м8\}4N����)��S�=��_Q�1��_>�ÐA�&\������8|3���=��,<�x5�y�a�_0Z��?���1_-��,��y I�^��i#�ɝ�B )��Q���W$��GԆ�J�G*�-��#�p,�1�0�2�������P]肦�y7�q�o�����~�S�����]q�,�w~�%�(c����9��Sr�=�����wN��I�F�2|�zT	T�,
�2�����՟Ƌ�x�1�����f��DbX�T�1:�%�6g%�L
m&�e�NŃ�v@�����^`���>�7jE���^�J� ��u��(EW�8P)�F؈�_z�VS^(]�'K[�B-��ӓ@�#������I�Hs��"U���(�����}9���,PI��}Ǉ��!������S"gw�}�ڒ��uk��;Q�t<�ڣ��E/����<x���bb��{O"1��"��a�*d��`T��d䖦�:P4��bû�+����!U^�����DR���k�o7������71�e�S�G����࿊�T7&�# ����ƴd%?�l���_������ٰy��܆hE�-MG**����Z���4�9Y, W����sQI>%�t)�UZ(���>�'ES��3j��n�i5�q)�r�wy?��΍���{&��^R�>ӭ�Z-�o�Y��7�i@��m={ј�N�e�Vz�_�|d.+m�c֖�s�FVjLt�}�����s+�~�8'W\Y̹�;��SA��o�6�R��I�5%
#U�L��
˃���tQ55��c]V���G���=�[�N�I}�j��n�\�ِ�/]����,���2o���q�A��������)m���!㳶�s�`,��U7�bl�{cǬ�*\i�����Fk���)x�-�3S�Ո� �����?�+�-7誵B�}@�=�W�G�\��7iRs�;\U]�6�C|^.�G��<#��Ćs1��V� �Z\A����3q����GXK�{�r �B���)����r�
�o��a�9�����x�	HIr���6	�T�������A����o@�ұt��[��8<<���<�5���^IuU!�Di!S�:����=�a{���Xebc1�y�ɖ5Z"H������">��?�䖥ϊt����)Q`צ7wf4G\�{T!y1���~��L��:tOD�����$�k8$͂��ȗ�T��]T{݇�,eI몙�CAd 4��21����29I �&�Tm�L�Xy^Oor`!�q@j��ï��z���7Jt��E����tςy�Ս4)79|��˩TH����M��!\t�@���z���/�W�
l���x���7�}p�A滼1\�g�"���#(����.�c��o��	QuT�uѠ6z����9{Tb�Cw�	��]h�F���:z����yBw42��ɁH�%gp���:��NY���;�-hg$��#�}42aA|S��O�b������M���Ɵ�ђn8
�jCs�z��TF�����\?Ӏa��_Ba�І9�_��JAc�Z(zN����	5o����G�7�_F|����q��?���A�g�1/B@�h�p�Q"�_� 8�Bv����F�=g�P' 쾴bm��﫛�r+�iR{��_�H!P��Ȕ�f�1��=Ӆ>6p�$
FZ 
��ddzT�}ॠW�@��s�U�Fq��%���4�)�&�J,5�e�������`���*
����w�<6m��ܤ�b����ݪ�n�*;d�{~|�V�D��?:�BF��!ւ���G������콣��>��WF�Re��� EM��2e�^����'y�o�a�O*V�s{���n��̜5����)�$���
����Rs��ZOe�&�{o��-���r/�F�E>�`jAk�z��N3�D�=�öKD�#\aH�z:�:0G���#M������q�}E& ~2r��C�h�7}�T�]ș�9���i����t#I�~Մ:u�(0�}q��&P��J��E:6]�v����L<>B�R�e]��zqV1o��߇N�<ƀ���R&e~��o/F�Jo������\��5u2�e|�ʳ&ig����v�6s��rs�{R�VrD�6^�8��(CBG2����H�� O����tSn�������s��͡�j�� Q�'�������Г'[Y�4�3Df��!��DӋ�6�H!H�K4o"�uM}�|u��#��L�Fм�&X����2}n_/+#`;��U��i�����w�]�֖��>�NE��"φ4�jqt�mN�D��?��!"��� �6V��3�p*�q׫�8�z�:�4ꛄ���C����6o�0���b�xI�4?�m�(�*Yz��Z�C���!N�E�޿��j�xQ��a�kҝ�̥�1!ۖ?>�|�����z��+7�ǣe0�-�߭z��{Z	 �U����C��OKM�
	8���/S����G��I V	\r�F@u}��ĈQӉC�/ύ� wI<19�V�NS�Ս���(�g�#z� �9c�sfp�V�b8�F������ߎv�u�j%�|��G���q516�[=>XF�$79���i&�͝�ؕ�ǒiW���������g��.�/]F����s������6!kw�7�p&{�(����ZQ�����G�ҟ��δ��q��t���W!��C�d�Uk�{:��n��܋e�ɵ�Tc���yrks}��~X�@��!��a�I�S��~��l5D�X�uA�>���C�ep�w��V� �� �7�S-qR�}0���E1G �z�D8�P����� �,���о��_m���W�����՝ȴl�������U�'�2��-t���j���t���B�ezp"���,��h�;���dI;��g��Q�B�'�x�ᄾz�tB�$m����_��u���H��!Ü�4�׵YRK�yAb)J�XGyo����F�æ�X�@m��6�\���#�e �,#��A1:�*dH���1)^����q�������v�hvQ �5��؋������T��"/6s}�|8̐��Z#w��i�˰4K\ߐ:։�;���m�e*ao.��R�{�I�ː�C=8��m�w��3<>���ޚ��{ti��k�%	�-�7�)/˗�����u�5����1̑cN��o+*g��^O��Pݝ��|��k�1���'��`�<�}�� �y�<{�])�{eBy��1a��Ѝ hf�r�t\hw�ֺ��EӓH�C��\j�0�>G��������ZI�{s[ki{%�D�>����qT�${�ɠ���'i���8�mL��{��=m���=�"\HZd��"����_��Y�>H�j(��D*��%��[������J�Y&U��?K���7x�\ۿ�ق�6���b9����J\#��-�^�5I!(�9	�s��n	�W����7gi�.f����b����ך|�n7.4L����5�C� c1yY�v�&n>��bH�u Y����KS��Ǳ�sc���5?�jZ����P�Qogg��1:)�b��5���2�T=s�G��N��h��2��vNM4��*����к��e�SN��o��89>�� CA���S.�����lV8_������YN@�����ڽ����f���ӞÜ���O�m���=^�~@vԭ
��b�;x�R��@��6+e�.���ڂ�C{�1屹�0�Ruݝt3�,�όK^q���s���b�s<�����PC��&6똇��/h��P�
�pBis�7������T��y����65@d�M��nܒٍS ��~����>A�R���7�vg3��≺"]t��$F�`ȅ"yH�eC
D������R1�Cz�+���e�A�!V����C�L�*��רLl�a��9�WQW�C�.V :5�u�P��$�]�iǄ	�l������B$�J�RB�m�^t����A $������oB�dxv\\i$w����7� ��j���
�x�[�VWXM�{Q�i2�q%`T`�X-�+����7�Ž}؎ vGFPP.�L���^�P:s�'&�A�@�f��M"�����²=I��~b)*o0�1��&�2J�	4@o�?���mbM��}TC�+��J�N����� ������\�%o�g�^I������Z�g��\>j)+�����GWIe�D�ޞ4�'f�E��
��K����XpP��|�u�T^@�+{i9�\����܏uCK��hxճ�_��^'L�m�o)�B��?2�`����ڐ*[/�$
%Z�3��t�r�z�����vǇ�QW�W��j����o�gE��>ִo���jJ�t�z]�T����D�^�dM��h 3CUiG�&B;CnjMĚ�c��I�D��yl���	<�#��`oP��R��L9���X`א�%7e:�3��_<��ԩ=�ܲH��@"�U��9�1������0b]���<{�Y��� Q�x�o��kD��[dK�r�Q��Xdl�k���z�`K3غ�i���f��n� �S��Z��s]����$wV��U���D���44�c�/��E��t7(m7�>D;�F�)�2X����gݰR��K9/��.�y�!J���~h�5R ��=S�����0	+�Шh�/�2@8
�3΅`��bI�p)"�������0�� �P��]�=��r��ѣ�+ҳ�U���1|{���T;<�0����,�m,Dt�~�w�'�Bm}�̏g��w�qi^e%�{V�W	����S2ckuu����d�7Ii']ڈ�F�˭�t~���&���Ě���m"�m��'㚀�h�
,�1$�lW�U���s���eS4Χ���Vu�|n�^����h�"t�l�lg��%HM�M��J��]+��'{\/z���w���	��d���s>$~���|&��=�,� fKM� �,vP�t�瘭���~��3�W
%��\�B�v��JJ/�։@I��cd��=�����B���Wu}g Q\eH�e��r���*u��o�hp��G㞖�Bw?|�&��B����8���x"7�b:!�p��!�C�v��3ȷ����&P�ʓ��5�^<̫p�(�S�;��a`V	h��$�r1�H�cݼ����e@��!]r՝Zz�m	���+:RPc����`��U�w:���0[c,�"ΓYh!�jA�����XO��W��$���h?��/L�;���hD��@��a+������X�q��֔@R���c֤x����Ɍ"W%~�hc�禐� ~r�O���OD��2��ʃw[�ύU�hR7f{N���G�Jǁ�x���m{~uNT���
��Z|��l���y:�y���׹����y�t�x��
W���}y�v/�#D��ς7N&�wIbl�̱(k��F��%R����d=L�\��7�5%^Zs���jQ��������-0�Q,qqzۣ.��E`_��O��\ԡ� H"6 m5aL��׋��~'C+��~]j���^�&^m�eC��
��F��@:!g�,�Mwf��H�<�`Ik{xȧpX��G��U2��,��¼Z���`�h�"�(�����fh!���f0���J`�X��;=�^<_U �y�<R�.Sb{B�
9�:d"g���"��d�wQ{-'ݎ:�����gq��F�z�yR#��-l/@V+�Z�*���Sc溗|]�*מ@�q���|Mh��<f�ήb徴�6ch(����}u\;�b^q�.ER�@>s���T�;��������3�x�e���G��7�1(��|.�3-ƶ��WBJ��z���)�Hg�ژݩbe^ȉ��uZ��zaZ�]�bW�&�����g�?X�6�55,����]LQ}�kl�\�8���p�c�@��V��8��m�S/I��,�����/�,���N�L�@@��Z"����+�T\+��@����jB�'a����{���(����%����j�>!�<LX�3�|�k�J�F9,�� ��O�#A��4{9�ܤSZ޿�J=[�`"Ȉ�dn��m9���(U$���2�@T�4��b�9O(/&��`�����rQ��Ac�C��Qg_��QD�=�m�f21$���`�~����p�b=T�s�yɸAD!>�
Lh��[��1p��(`�:t�e�y3ڛz��>#~0�f�<�)�l�+x�/��NyPX��l ��o" x�/�T���Cߢcsg�T���x<�&d��tcch]��xn��w�l��k����|�RH��ҏ�
ę���p�x�q�H�J{&�@��!��>Ln��{� o�h�x��N���F��-{�W�t�m�fN��{�Y�	|�D'X�kK	��%�`B	��x��-c�v��@��O�V�J&���m4�:X�/�x�v0g��J�J&φ��c�mC´Q;�O��e1�f�L����w?E��S@�,x�k��S�Uk��.�X������-s�'�>�'M�k:��]@���ۂ�����Ĕ�
�?s�����W��Xo�Bؑ;ҔeCB���Z�[d\$�ng�F�W�-rU�s��`pCg� )8W|�-�F�,��Y�H�q<����4���*��C��p)1W)�N�m�?ݷ�+�����ĩ� �N�y蜱�j=-m�FTg*<���o]$=w�|��sf�-�"�@����L��H�ͨN�}��[�p޴������4*|��+E�{Ȟ�"�[���o3A��
�3J]�L������GO��D=���a�<��.��ۃ/�"/!k��ۉ!L��-��U�Q���D=��8�\%���DZ����Q/�T?,
�N($�Z��wl36Ő�K��� �c�נ�9x�0P �����pX[��-	$��$���=:Go�������(w�����4-ԙY����:����)�d���2�x��j�/g �E���g2�6*! ��N��E�IIEG>K�U>H��|L����ԟL����o��?`�9��-7ua%�Z�ά��3}\���,.(�vOἍ9�61�JC�0\ik� ,ŌPA�o�ɸ�UGf���-@Y{[*�T6Lϼ#�[��h��#���F�5�%�E|�^"%1(�4<�SV����P��3�q昮Ԑk'D�!�5����K`�E�ҢL�S�Z!����#��.Ge�ʹ�s�&է���$��������O�@���,F��7]������9� (�e�in��n���/���L�Z��q)�?�lsHsw#�����j���t1�I#�?y�v%ޭt}����JN�e�E��Z����:A?Pus��C	��~�v����h�p]a�� �L�ݯԹ���Υ(_��fC^py�l'�,9���D��KV����5M���#9Ѧ��,hoǆa��Kh9L��tii]����([�0�2�)-�I\�E0 ��U�yڼH�e}މ~_7S[h����	!�b-=w�ee��)��4�:B�����ev]�F�:le��^�Q����NcWtE��I����& ַ{�9?��x�#"���;��M�$�Q����ڝ������[6�L�=��EY�^�4\�f�����V��7�������7�A���*^�HA�� ���aG���5,�	�I/�5�᝟?=� �Tq��L=x��C�@ޒ�tf�b�I�֛Y�=9p�s3����^@&���M���1V������Hz�cC���L4��A֙���^>T9H���2,�z'|D����!����G@[t�!��F�C*`�B��,+)Z�/����#����&&&����b}������&�	P��߸�����	�.��B��hA��-���y��k�졵iX3�������W�x�A��6̸��(^�y����r`.���\�5�����Az{�Q4��|�+<M:�!8	�Y��)���+W��dn�Z-�p���<����C��(�c�H(�d!���&w�hh���T�Ⱦ��q��F����F�;�wtpř(��)e�E(&t(�9AHK�7�yS��./�$*� *� �O:��7PU�'���P����u_,P2�ҹi����G<���� }
l}�����V������D����V��ED�����~�y['>2uC�|?#?��I\٣�(���-��1����P7b�\��l/~����g�[�{����]%b��lUE&�`{W����x�?��g;W�9�?��os�:L���?�~%O�E,n)`�� �A�"�y�P�T������7�����7�fI���6����f$r���T�ҽ�[�/���]e�&p�E���ޤ��l4B©iD�t�ўO�m�B^T�V��e����!�/���|� ����e�VNT������׳������V��c�`�M ]�nl`i�?��wN�a��#�z 0����P�Yw����&��ͨ}��)i�K{���'
��y�#�5��F��B��ߣw&��Z���|O��<��`���mA��ҩ{����7;uN��/��L��-Cm2�  �q�[4�Ӝ�h�m�PѸ�l�ncov�*Rt]�Rq��
���V��ē�L$e��s)�*}0lK@�==�)G+���&�xM�����-tgqr�� �g�$�v�ɩoa�oI��V2mJ�$J�����L,;#R�X�˱�~mD�r��0�&D����B����� j"�8������B��R�`�߸��� ko~��cF4�g5' ��=Po|���V��9��B�{k��n�t�0QK�IZ�o�OW{n�:�����Di���y��W���&�I$=I�k5��n'�Ei< ��3���\��H�b��� �����<��`�o
�p�}��棫���ڀS��KŘ����P���tÛ��C�~W:Qό�C<����&�<���d�K�n(�V��v�AE�� �:��j5Y0Ӡ�^�Z�!d2�=ev���ų�%S�6�Ѽ���LO�V&��oZi��"�Y��Z�|��v�,rA�JG���[�AP�fD�M,ZeU*�9�b�E8��^궴!�|�Es*ڴ�t�I�V!"m��X��Ĭ�Ǎz�cx�;¥�c������z�3o���"
��~b&�#D9~.��0�����'f�� ^�D�����[��3_�7Y<���͔2+~g�4�/i�)�S�m�HJ���.��q�f�U����5n��\%-���znb�A���	ўr�;6r7����~O�j�}e�⬞d��ٶ���tB�0�V!zgF���1�Z��3^rJC����T�p����p�=O�nT2����=q������k��������5ѿy*j�:u�6��\��oKڪ���_�3~ۯw�BL�e���3!�,qwƎ���9顄>P�v&o���cܻ�� �ADB/AA���yl����@ҋV�$,��I��cwW}�ݥ�%|'FY��&��u��׋/�w�mp�7O�
!��aK�4bF��rC��R��<�^���C��[��T��`Y�ܪ�i��T%�%3pe�9�R.���{4X|�_����.v�m�a�y�V��C��Hi����E=��\Q+xZ� U�ԛ`�ԡ9����y�IAW��Ӌ,���G~�V�:t.���I�g�*ОK��;�r�z�����,�b�yX��+<�֯�[F�r��=��ݶ��D����`ΩËnjT?�b���L\YX��Nr<B,���.����� ��C�}�|}�$0��������-������_Dh߲�����2�g�2
W���L��aN�����2$`�(MƧ�]7�xh����&v(ၬ�==��2�4!��Th���<Hģ˭.���M�����X`�/��#�3*����F��;UL�i��%
�o<��-�nTj
J�rn|~�����갩yQ�(.�d`,���\�*+�0������C�s�˳Л�u�9�H�4��.9�DP�q���Zp����D�Q��=��_
�ԩ�0c����N�;j4 �Y����Ϟ�aP��q�s�rjR��-�����+z3[p�y��SI�z?�|���y0���%���"5�g�ə���@/��S�ic=G ����D�xĒ)��5Kd�d�K&�&U��5Lp���b���W�F�S�sZ���I�e֔{�� ,vvQ�	�$&k�}��o:�3�y�41�O��F)j�ya�֙t�
�0�l������N�_Lv���߅�o��^��;bD��wU/���������� �u���D���W��|��:���
�O����b*E�-;>L���I��W�c��Y����AM�g����l�G���� �q�Ei�5���������������|X�޸Jƴh,ʔ�w���f�U��4�#k_	�O�QĔ��PU�w�?_6�����%2@��5t����!\-R,cH~M\�M��b�e+:�w`݃ү#TCh�]]p��&�Syil�^��+��f�j�6r��c��ܶv���T��1�qeoCxY������<�E�������סW�l�8`(���J&ٹ�a��kkf4�C|��Q�]_�x�K���b�զH�9�b�rv߀�Ѽ����!.��9V�̑:�S�>o3;n���Z	}��H�&a��Aq����T듽����,��E�)1���;Ǜ�GB�](��B����]��|���F����F�V���Rq/4]��]n��?ў��ɒ��h��=&���=Wk���x���K�(l�ӭWx�6(����|Jp�}�.��*=G�7(�i���gN�O� �P��,9����m<;Q������mQ�����ٰ_����+K�"��a&�}S`�I�֟����6��e�����[3�BD<�q&�2l����i�F��AK���`#�=�R׋��O�\���C�e�K{ŉ�RZ������D�t�2,��[˨�>�Y/'�mx���'R���l�U���	�A�#Dax�LЁ��y;��μ|���X��~R��� ��o1P\�|��u�^���pa�ߧ�!A�X^���<TV�x�d�� �׆z��sJϿ�yh���e�f���^��,�����Vp!�����m��/�a��d�X���"���:�	;rኮw���m��a�מ�c
����/�)t��?�#n���v���q[4p�>0M5��<���8���`ةn�s��D���X7�2o�RsxM����MεD�6*���Ѯ|����|!�l^?��j�a".o6z2�8$@�fa_���<����[��`�� ~�?@��!�� 8uy0!��c�v纅� M�c�`9ݲ����R�#�s0�1�$͆� �}�}� ����yaV$�A󸖣�݊j�����4B����$��$:��0��q�9�PG�+�ɵ��V������̚B!�q@��)� c�X�%��-�dg���M����W�:�ltJ��T.�ZugFmg�e��9.@��K��V^*��8����4���:��)������J�8lȨ�Z�ٍn���ғ�2yJ�y�+�� �,~���8��?������� ;�m�,�P):�
K�Fۮ�`C)@�h��gŶ�X��2���S�8�3Y�̃p��MT��m��gs0	1V�zI)!l���G���
����mU4תa�79V	�&�tQ>�Pd}�p*\�?�Ɍ���hDf�}-W���ԭ3��vA��0ϰ�F�+N";� ��D�I�κ�ui;~Y~��C�׍�*}<%$cY���o����+}��~u/�PaA�uD�k᧒K�`�Y��̨B�^͚�{}�9x#Sp���9�k,.}5��O����w��>���*b����7bC����y>t9���N��ل/9��"'��@hR��A�u�[6��Ā��P��W�#&`��l���Z]~ �_l�����;8#�ga�����Ng:���s�����A�J�	k��Q�ٜ@/;�Q���F,�E�;w� �{9�՜~���҈�G#�J��e�=��%����J84 �<m=���ڨ��%D�#VI�s�}�Ա�aA�*�׺ul���%3��s�/���~"�V'
�V��q*�ʌ]��󩻕��{���ߩ3֒�i��i�Li1(�^��7���q��"��p�d�fkԅ��6򕛷.��;̦Sh���	�u�(w�A�T�ʗ�Am�+�8sfT؁�-nXw�I�ռ���mbok�k34�<�p��܇7k4[Wc��P�{9y��J3��.��A��SyeXN�b�CzۮHH`}�����^ң8�%xt�e�mI*��&R~��6��^�ߋB"g��H��	cVQ��q��o���ߵ��������5EgP"\���O�j�o�#�L�a�)G��zZX\v��1��D�`�a:fV8�l�J�ln�$��p�$��Aj<y��l����d�n0l�����BTB�$��{��R�P�i;�#4H�F߁P���1E���y��m�y����댱�����`�ݿ�r��`2pu��m��q�խ�[��~tg&:~0O(0;��j����'QC�:��
�ʔK�6��"�Jxxj��l1~���VȻ��;���UT)g��(����Φׄ8 ��8Űqx9s���M�O�.������W���p�C���x�e<=��j��Ϭ.r���:H�w��I2Ů�Dg� ����s��6��}�/_9$f~a�,�KG"�F�$�	��*�N�| Ռ��{�9`�b��R�P�g�FM�b�G�lTcH�PQ��7p�-��	y4��:�v�b�6c��q+\k�Z`G^?�g<�]�����_f0��eW��� �v�Ę���Ni(��E:l�d�X�G��[$����-�?��	�Ci��Ԡ���:�����u��Q�7@Q��2M�X�v/�;G<��+�M����s�=�c�6� {�%�Q��������2ч1ǟ' ��v�T�4��	ggl��N
�%�Y-��(Ov�W�,�_d�O�fc�2>���F]y�O[$�`����>�o$���d�j�+�}}O˳�RG��t�g}������Q�	�7S8J��o�M������iѮ�8��0�ӒՂ���;A�ڏ:�)�Yz]U?��w�ޥ?�_i+մ����O�^o�9_RY�����i�fNo����B���xǵ��`�4�:�?Q��7� N�	�"�75���{z,����N(.S����ipd�/�F�cQ���}2$f�G�F#`����"�IҾ�Q��rY�ft��e0����'�W�|`+��\'��EB�=��'Щ3	Ł͑N��L���#��xk,Gg
�JW��Eem�p-S���c��]�������?]D����(CQ)��嬥�A4Г:���,9�6���G�!2
S�a��O������4)t�>)-�	~�ȝ��v����Y��P�?�$���@b ��D��[�
�ߪ3zf��Qj�u����!1L�\N��3��Қu�@��y��:���؆�q��U���l��͋Om��=&���l�����aAV��+W'<_�$���Avh��UN��)}߄7J�O����z^wmc
V	T*NA��~��E���
�����Vy��	p�1�*}�����Ǝ��`ꕻT������ �A�g[i�\��?���H6�. ���h-�X�h�7K� �2��Z�=�q\~O�=��% �}P�Ԑ5om�tRH�A+=]� �Ju������f�{��elw�hOc��r\˻�)����1%��=I�޶�Rv��֒�8 Xg��y���x�ͮ���F�F&J����Z��_�s���/- uP@	6I����I?��+v^��E�[僅��o(�t�(�jY�9��Q�o�^��7
%K�@M�\�7�絨>�s�W�
��/����fG]`��N&���Vē){�c� �g���5[�sXx
䥽O)�X�BL��`ɡ��TJ{_�`�د�������'pL�)��8� ���n��-�[H��\za��o�8�,�7}�pN�����ꫤ��"!Y�|I��7��Xi3�VkD��e���Wŋ�4tvr�L`B��{`�QIX^��B
���r�Ejv��T�);zV�̈́���Te�[j�P�U�����x��S4��HY��P����� ŵ!mN�A��w�.�@��Oq�W��o�aU26Ty�+ԗ֔Ĥ���ȷ�$lhw'�6��mٲK�OU��>_@`5��*���gJF���b2^�k��q�m|V�3"�.I�lw.q����#�SG���k*E-ph����6�2!&z�m���ݍ�E�]�L녫C��4��ı8��U�O�����Ў�+>!��.q�/�wȍ}��/�šZ�:��[tu��(�q��|�=�����Aw������ph-��;}dFG6HL@  =�̛7��w��~[w5;d̯�n"�ȫ���9�/� �jA���u���A"ؘ"m�dG=��˜dR�FhN��W>�x
/L��JK�S��ߋ&7Ǔ��a�Ӡ�n���^L0A� ,	�p�����C��"؝}��=���h� s����y��� S�v8�Vx%1f��Bܗ)-���2x�@H��F?�!sS�Q�0�~X�`�}�LU6��=��1ڙ�>HI�C�:q�H�(K6�!�k�[�-.1Kt���U��k�L;�ŲU�%�T�3�T����P(yD*urw7rB����{~A�Mh6T?���^�V
ǩ�Ra��ݣ��1��Ʉ��9v�&Z��H��v��_�FX.]�Bj壦ͤ�B�ms�5�2�IW�rG9J 
e﹖';)�sY%��bs2j�`�?ؓs �ܡ�W����Xk@�ZN�^�x����GBRP5sj�e���
��֐����Yc�+E��Q>ûny+aGj��Dp�z���#�,.�A��nj���3K�[|��pF�������XCN�=��&��PZ���t9�е&(�3��ݤꇡ�`�����K?���ǺЖ��i�c�#�<�s+� �����Yv���0\��θ�����Zs���,x��g�6F)W��[�|�8�r�.=����܎O�<�����ELyA
9c+x������"�4,�
���uLCI'�0vh���?�}�V�7ST�jŹ&t	�9	��.���w���93 wG��n����:g�?�=��G{Ē�RVL2{�,���]j�����e�%-�Y���°��^Z#�<�*�Vޖ�#
���S��9X�ɥ�\22E�"n"l���ҧ���i^��'��v_;���f� ���៮���3����L Z�t��/Aĸ����[߼-��߄��`ã�wEn�\����v���R(?~�#��(/��9�_;[���SO�IѶ����)걑K���G���>�~T��܅��lf����������#^�vn_�I���\���3Ŧ�q���{T���d�ɏ�|a�fX��u��,�)K��J�vSD�v}�`Y�b!��Յ&Z�Y �o��W,����o�0F��Y���Yuڣ��� U��E�3��̐�e#�B�h��*\��o�8)�&�9h���P�<,q֭V̼��˛c%���Ӂ�
7�m���=�R��=d���iMf�?O�al��q���0���XU�t��c��_�� Ru�m8�M�E�ϪkLb���h��Df�[c4̀���6�Ē�'��4��9�!�f$ұ��VqtU�O
4J�m,����JU��Ց���p�Pir�D؍�l��)!]���P��}wkc��t�f�s#����T�1����V����-z����Co��9�Ϯ����"��J�:��F�T��)T�~��e�YDK�bI��X�f{
�;mXlKn������G};P�3�7L�7�w1[��-ӴJ-�3�S�Y�hB|�_���
�zl�|����&g�E65�`�G��%��	[f�	�Z���w��.Y��r�>a�#��4 g�"7�BO������;#���Y�������Y���q���<��oH�����vb�e��]�,���7R���H����A�}��B�!L��>Q|�pV��$���KFӻ]I�H�|.'QY���H:EC�%�B�u�m6��E��A�{��ʗ��'��3��(���S"�_�k�Ѽ���g&P]ř�0	Ԕ~�ʇ�Z�s��|�]���|B�	m��f�3��[=�	8ޘ��Xۋ�N�ʳ��~�mR�1��=��z�=W���=z3D��o������
�kA����{�*�h���S���@� C�2��y��ݫRJ�+ю�Є�Y����嫰��"V�@n%�	ʼ�T[�jS���U�]#���%�z����Ƭ̲\a�z%��y��T�[�Y$�JD	#��7HJpGy��$[��L�4Z���/�M�a����<����,H�^��FN*��.���=rmk;�;��.���PqZ����ƴ�B��%>�~x��Z "cX_]����y:W RF$ՒF���ހ!�vz�9X1�_��ŧw�˟!v AZ'5�/�ރ/�l������U�O�޷Pwq�@�}➆%����Nc�ϕ��>��r���Q͎���^g��.KFȺ�2���2��r�U�+e֊uSy)o:�����''ԉŪ�x�~��r-�.D4<�v��H2�֙�̿�u(��:��a�$~�},Ʃ����Ǹ(�
�]��V9c������Qߥ��7��]K0T'�RXU�=I&�C�Ԭ��jVޔ�@�M��1dn�k���/��`�����1cIU���0Þ���B�fJ����}�~�aR�|�G3 fqq'���h�;�^�t%*	��--�.�s�����'��8�[6���Su�#�����?�_:�B�z���zOu���%�O���eԄA��W?�1��sj}6m�]ATZuDi�Sl�$���gC�q���l7�bd�����@
f��[ɠ/t/q��$Nh������`�(;�#��d�	 �u�p�	H��KLa�kk�،�K�^�V����q+*�2�s?��+I�=
I
 �
�Yf�THĨ����������9�	�ic�o�T��M���:XWL��Y�шg*��A�|B��1 I+?��p3\���p ��C5�`�%�R����B��_A�ĩ��{ �!���~�K���cx��#~i`3�bFtJen@<�P ����Q�� /"����6��~�+�h�b���v�?���?�q�%;\,��Ya��?C]TSKW!2��]v^��<=!AI5Y�gr# D�hIϩ�v�� ������8s���A�.m�S�O�Q���?�}Riqυ�l��k��uj�`V_��{qH�H'ǂ��KK@l��'t�a'r���y�Aܲ�#�9�ۊ��'*;C���X� /���L�u�ϛ��)�@��(��	|̱}-q,4�RJ/Ǆ�-�ܐ*1v�P{���Z��톊�j.���/D^��l>��2ȓ�\���e�a7IHx���j�����Z_�te	���G�V�_��Z�qi� ˊ�Bb�;��J���h�(�������?�A߶��"���:��x�[�o�f�7�l�d[حf����BR�*���ع�_�~���#�ۆ J�h� �olk��>A'�}1�K�ϊkW�W|jى��}�1D�bj_�|Pt-��j�  �_�X��_J1��B���ҡ*�g�� ���i�b�>Ҁ��rXgﳖ8��&7����*�/@@Te@���6B|���R�	���3n�G#T�_���Ic��g�MN��)�\N��4�:�8�#�G6W�5�7��ޘ�)�l����~���&{u�i�������vH ���%�y}�;�c�%��}�*�ݴ���<�\�Pk!x�_�)*O���I�(�"P�GvjD����h�q*���m}��Ɉ���sQ�`;yNڎ�{��Ǜ��f�tT�t�A��,��2�e$��t���!�`>P��/2�#{/�q3�k�^��/AvO}��9�"]�&��[�_�J����.�/�m�V[Fn�$v���̿���w��IX��7�>��̚��\0���(j
ݲ���� �,�D���ݲjS�:�<a2
�I��k'v�K���Z:� �
����l�� \ݮ����������c�g����L_��(�J����.���%��E5Zvb����bJ�Jì-[PS���X�,�8uR��Ş�C�u�,Iny3N�c�'f@���Cv�Bt��Z������cU9�4Ol=M~zh!N�[��ۤ�{��:zS(��;"B��wg�:23}*�M�oj͗� Q�����Q����Or�5gr.��/�."�x)�D	���2�����x6 �`T�	��~�����3���M��ݐϼ�Xh�������sgfk�vG�ϑ�����s�i��6��D�g�����<����XvoU�/�ñ����{]Xs����r5�@������oŢu�z�H��Y=�
{DK�5�LV���C����E3P�ʠҔ(!��~��{Xy�@ag��7�ܰ�S�m����V�u5��� ��͎(���{s�5l��f��25L���*-1�['��ܞ���C��d`��4ͺ%��l�#��:f�w8j��k���3��J	���Ag��}ڙ+�} ;,�~���3���!��E�[��&������𸍅��B3�f��[��z�O�j/�Y��B���{�yR��{�����o,�y#��lz*��������h�~��z{�FO��Ħz��ڤ��T��SS0,n|R�Pa�A��q���+*y��f�B8UMA��`�@"�����\��0"N����=t��z=��-hĨ|��l��H5�=�q��|��2R��HS���R��cƮ�L��B�v5gK��~��n��$�m�ٯ��ci5��c�(0���l��� �54^']���ebح
�@�mL�3��Y��0�p@�y�L"# �`F�ܜa����,(o�Ʀ�`O�"���Ӌ{�Z����cr�W�[S5\$O1ZE-C{�C�� k�~	�:�*W��6�,�f���Nf
MB��v�Xyx�n؃��Pdx"��bm^�2I�ʅ������6��z�.Zҁ���WXU�>'�)Ec���f�~0�R�Yw�I�ۇ;���CR��f�����o����1_ �R�H.:��VY������>`w2��#㣽���O
��q�NW@S��9�Kg�G�KK@F��P@�e�YNmL+�a�8�|�%\o���!	��jr�j�ؑ�V7��-d���9r��3��>*��wPq�,�D�	[B�V)�32���*��]Xӥ��<�Ňqÿ>�(Y�72�l���,�h�����ƈ\�<�2�,�4]����
��Bꗖy�[k�#Wب���-ѦҶ�	56�0h��9ĵ�6�Ԓ�i�Xƀ*h폗��㇣��Z�
$����61*Z������*���L��i��=a��+�wp��l�@��;�3������Q+���P#p�帖r��r��0�	�),�3nmԝd��sg�U�����]f�� |{!K#W��>^k8�����P�W0@�]E���K��z"��b��_�M�8�� �o�����aZ�����r{�⬨d͗�	T�c����Y�'6��Duϴ�e� �Zz&� �2�1x^�b�C*�3�/���'�ì�Y�BZ�d���n�Va$�^<>tO�/�?`fwL�U��9>�^��W�����׋w�2����9�u�?L�-��S-`�<C7�P�<)�5hDۃ�;�`}[J�l2��8�y���ߌi�@�
��".���b�s�>���)ؖ��<���1�)��Ic���F�{�f�;gUy��L�'���]ƫ~k�VX�EO]��է���[C�E��唱D#�qn[aev�v��V�y�����ys�ۆ�%O��%�o%�+?�+MFO斋�^�G�˘dx��[����T��1�9qt�*�8 '�lZ˙�RWh�=������X==R��LbwpX'u0��ų3�%��{��'���Ⱥ_'�����)��G�C��D(a��6/�A �.L�@o%c��y��B�N��)k�*��w6�2Vs���Qs���b[�K�M�OH�lTf�ۆ���x`�9����r1!|7�Ƥ�A�~։
�e�P8������+��Q���{SA&ƭCJ(-Z5H;�qx��8C����B�#�f��� ^LZ��3v(�A��}��ݞ���ѣ�{�9!��%0����P��Ƈ�/�<����j��v�}�А�5:G4��į��lȝ8#`�į�*�I�^6�^ �[o���sT+P��˩wEmb8d���PA�q��ی[�}�����.b��%/8�Q�M���9��ʘz�	�0F~�=�6�n�?H���j�-��$�	BbR�ε���upcC-C-�Q���<
�� �J3���[��.�m�Ͼiz�Nx�6��~ۋ�l}gmD�$�U�]͟�J�\��b�)o�:�Dx��>E�z"kLZ�nх�����7a���ɘ�=X\�3��<�z��@���*�Pܓ�q�!}*i2MZ��������N�-IB+?��$��'1>$ğ��NG��a;/����A�yZi�ȿ��X1�걶`�>���lnZ�@$���X�@�!M��,$�����G0k�7���]/&�by�Cnw!ty��|KnX~%܉Vc�}�t��Õ�3���H�L����2C�s�z)Z�z�@���
�]_��Αm��*1~�kJi���qK�)�k?�4z��H~�{O��5�f�p/yT�[��;=>�>[���U���������X�ѱ�-U�����-MB%�Vzx��~�>ܿD>�Uݍ��]U#����iiғfIǜ?c}��
�)2�w	�d83��R��Ԓ�!�«�D3�O� ~�Q�VB��-K�2�},#���ǢJ�5��Y��"�l�u-��'�.ov����1��4�u����~?�AF���b��=w*��w��3�f���� "��|{�������Z��$0\R�f̴cb�����{��_�Nca��]2����3٣h�#U��е��Q#������N� �*�،�6��? �;�6�tlEzr�::/z(G��)�-JR�T�JJ�o/:��7�[��K���a��A'ҮV.O���P!?Y���|���I4�A���U`�bw�9�\��2Hz�6|�%�%�Wc%:�]��BM���'�$�/���"T�$�2ߪD}M��R�a�� E�|��\nn�$Ӧ��%�:�Mea{5�d�Bg� QJ�8���!�bQ阊Ċ����WX� 	��b�xY�zLM-�f��P0�
�SNN5>��O�䕔���'M1����I���yð<�V0�y��G�[&��,�ߣ�j���X�K��k�0�2�t�)���ND�9t�2N�[g�V̖�E��=Ur׏�K������=UX
�E���t~��\"�b�����%&�#�����ڌ�dR��%���||��-ۆœiVoz7�`^��PM��#bD�#ݒ��-�/��;Nj��4��i�v��U�E;j�򭶕T�9> ��+=���kS�6��+�¦S)��lJ��{t�=�_N��� ��ɷ� �!D��u楎�.���: C������z�vRx[gv�A]zo�f�hL}����*;h��h6$фv�H]N��o���,�5�ʕQ���)�XR�8�j�5d���0�<������܋��g��'�*&�%��{A��I�ۛ�@���&�C��p��k��)���,J�L`�!���SVlV�̥��j�(�s覚��̸q�����w���`)��>H$�2V���)>y�����w������D��3��;,{�J�I�����n�-���$Vr#��9���JX�#]ۦI�4�:�ܗ�bSD?"���h���]� ��l/`P��'�* ��_)A΂� .G[�Q�O�G��(��%��*fl"�=AMצI#2^����:���	��I����a+Zv%�Iy&�#5:�g<�/�[�ߨf���uœ4�H��2��{�f�>���q|�kB�/{���p߶U1�.h�bΉfV�.
�q�^я}V�u���#��Xaq�c��X���Z)i|5no�zRc� �XdE�
r��E���HȌSL��bF���e����Vg�:��7oO�f�?�\�mqT�-�+ȇ񌘳k��;��ÙcH?�����ۊЊ�f\t�,q]�������A���	;
�Q��UP�ƶ8e9�aP�)mV���W��<�9��!�Ç.GmLgZ%�F���I4uxzoD��3j�G�H���g�>�3���9���-����"��c7]kXy�V:N�N���#��^d><ؒ�dx���[c��D��@VsyC�
$B��S�B}9��Kp�\�(H/W�e,���O�'`E��;�������z�$]�MH됳B$�bj�ӧx¬�-� w�a�b�z8;t�	���KV�K�t�r��[�@�����:�xXm�b�1��䋔Ѣ��B!�p֥q=�)v�}h�h�Y�i�)�nM��{��!��t�"�₶됸RE� Z| z��j�D� �O�u�S\�W��o����N�/n�z�g�8�(���I�ؖ���#�H�m4��C[��)sR�|�|?1L�j�Zy��R
�W|����ο��:z��QiE�p||�����E�~���Â(��1L�����53�� [vQ9�+IB��<���(��-���b%Q�����tG�v)����2��e�8sF��!���#��jm���
[��?���Z���v�v�)��@�K^�a�3���sJc�j��rj"#|���u�h��I��Ѕ��#���hEJAW�>���t【ʘ��3!��"���x3���<��~6{�|��J]������ժ��]�R'�o8h�LO�B� l8�����������3�׫��2�3����[*
�pXa*��k��b%ff8�k��^1�h9q��]����b��W���#i�6�����+uz�g�������g���<f�Z�0�{�ݷo��7�/��J: 7��Ǒl�Գ!𝀞J{D�;���0�h�w`��%uT���~q���PNb�*��r�B��ܹ�s#2�k>��<�&� �=��������	�#/2�C�l���C����w\$RV�k�Ӊ���u���i���#�[��	Zo	�pN��D0
�?�F�*H��c���,ڋyQgT��Q��L@���2��3�K������0}H{͈!(	D�ٸ��c�F��o�v��g8i�=��V@sV�UO��!}��$}U��S�[��M�nxE�X�S�E)�R]=6��"�7�I�dt��}�!
�
+!Y��J��߫:�q�2�o�@��
m9*tF�Z@�h�6����i3(^=7M-��In��B�}�&6�iq�y��%���e�`��ޘy}�����j�f&E7l,��4�����ؗBq��ŏa��\i���0�ܝ`đh�m)����+++�iBr�e�ѯ7��E����B�c!�=�XN�}8�E�?��^��u>�AB}<�;�G&�/�k,78�}g�>O~�G�B�&�~��wȪ�q��9]�+�Q�P����p��]��g�-�N�&;Ny!I�L�����w)5�q'Tm�x�PX�L���K��x0�8b;���,!����U7�Z1��ܽ�Fo[�^G���ͻ��%&��ě= ��%̴�6`���Om7��a��ֺ���O����Ǚ�;��B0v����V��@@���pz�(I`s4JP�*qH�-MK�C	�����(�/�"��@��*�Ms�9)E�C%�$�Ar#�g�Mm�&���H؞Ɗ�t�L~�>�	�*�Q�;"8n�ؒ�����"�}�5l��Q�˵��|.n�%��+ARP�\��τ,|ӑ���"5����9�	
X ���F�w�����8�o�rˊE�ꈼbFN���*�t��'��o�1����P�Vɕ����BB�Y^��6�}�'��{��֮s\�����Puӯ��X�I��&�c�ӻ�~q�+��}l��M�����@9&�}N���u��oZռ�K����-�@����0��=8�HTd)�°p�Ѳ��dLM�4�ˈ�G������w#�S~vr_C�Qh���Z�6+D�")�1!]�7~�l�✈	pbo�2�*'}��'#��J�>� ��f[C ���]e���E/�N�0r6�eB�)���"�(0�����Y�!�-4Qίm%�� �w�D��]f�_���_m� ���X��8�y�gdx��U �!�j���a!��^�*j:��8��^9���F5���kem�8B�%K=��s����x�]4��H��?��>���.;k����>�j��	�(��K�;)o�/����9��]�X�v�a���[i`e6C��O?<h��^���mhB��cY�>xb���:���-��ܛ��!0�j��W��J1��44�{�֥gS�Cz�d�u<x��t���-�2��S,j�T���oZ�p�����dG�,7�LU�N��ϝ�H�����[G���ٹ�e�F�j���4��Y&�v�aZ�
>-˪�m}���ʷ�+��ɏw�M��.e�QmulKza2<n��0�)'��	:1�T��	�O�.��8^2G���Fs�K`�|���X����;�(��\�-v��u�c皟�f����W�צ��,��_y�?"7�_Z���~�"^	�͡X��LI���� @1����ӞL��0����Ri8�ŜŽ+��#��MM����M����~"l{;F��<���=���gK�s�ڻ��+�������QP_|kX0��X�Z��2t� �g\o��x���L����<�w�7�t��Էҷ'c=F
�7����>l;�f�����8{���Y��-5��g��P�c-B8�2�D�������#�Ulbv��ɷ��Rn|�s�V���N�5d���~+b�)���<�)���h��>V��������҃��Zhݬ���Y~7)�^z�:����&:B-���l%:�oD,�{�ĳ`�V�1���5��h����x���e@���p�y�9��7C�?O� Pawp:��?���(�C�)�M�j/��^���/�;����} :D�(��Jm��0�O:DRAh3թW�����܉ٺ�U��f�Z�o��y�Q<����.q>�U�e /�g7��݉��f�1��p=�6���W�ם�TnH/��MB�0�`

0(��å�-��z��c�h�Ì1��Zsn�b�Y�n3�g��6�tB��y~�y����Q�������f胴�֌�)�sFy��S �K'��������ӵ{�P�z@ϏV���g�`u��}�XM��t�����9h�2�z��A#��V$�]]�4�z�;�8�{m��\8E��t��E#Q6nw�^FVMt��_W�ӌp�����~f]tU${��ˬ���������nՆ� B��V��"L��}�a� 9#,�	mhb���� AX'�{�-M=����J��l��Cc��������H��q76H��#}�8��K�!��7����_��Rڔ�*����u�`�(��VeS���6���bGU������F�S̦Dg��]�a�Ar`[�.�yt��9��p���zӈ�`�H���i�[e��.Qc¿���E��h�	�Ɣ�g�ƘL�(��١i϶�zV+�z��g3H�	�7����cy/XJ��ŕIǬH��Z���i�`?�YlVԔk*��x������4>� �v��;��t"dV��E�¼wĒ�5x܉~���qG�U���*c[nI�(.�	P _�����e��IS<��CH�PJ�MH�d����O1|�<8�A�,_$�oE��K��B�/酚O���� ō Ma�)�)e�ߧ#��3a�3Y~��\��%�z�zՋ{��^VU-�v(����<�o��U���I�w��DĮ��sD1p��N���@_���Ih�/v�����%&������ѐ���a���7�u�t3p�1P"D~yik���"�x/C!�'v�P�,!�uF|�U���i�R9-)��E< >|S��k憜ٻnoY�W�b�|K���u�fk΀~�����l�r�Ղs���ݥ8�>�� �E���F�����+JSh�#n�m4��P�&i)F��h�u!�.�Y����'[�����O�H0�3k����Q�sLPr��n>!Γtmť�;�����(��d�GS��AE�Z�@�L�?2�U�<�de%�I%}>C�У���\���r��^�x	|��}X7�8f��yp��9<SϣjF�+�C-KK�Tt+�)C-xF���I~�ލ6����,؊c�@a烆���)G�BxMl�tC'
2��g�s�M���_�S�U��Scrf	��"�Ѝ��/�O�x���o��Eb�)F�ͽM�KAixl�t�)�7S����t�jణ��*���P���?�Ϡ8��`P��i՟S�!+�b�_��F�@��A���:����3#z%�Z����=ЬP�	P�9���7��Ė��aY���/�>\	�tH$���<T��>	4\��y�Y$�<x����d��Ts��[zH�w��5�|�8��� ����H欃K�kb����y��E����������k"�ȕ�C,�S��6����ƒ$�(�0�x	�Ĝ:O^#8�a/e�׵V�,A�en��A���A��&,�V�pH�T��ڊ,�n=���C>�ZY�L�y��5��ޟW�<lx�KT�&�����0il�eG���iU��*���>�0|
�c��z���
�S��m�%F(Ȟ�اL^���Մ���f�O�j��iP��K����'©�_�Vk�'�LQ��݆�L���	��OW��I��#Xz�]O;���.#�4�?����L@�?�	cb0.��
 ���C��
�pLXٞ��7�Ӽ����4�_FI��3-m* �=n����ڒb�����3f��z�.�z����G���Ѳ���9Csm6 Iho�8�]�+�:�I�3���/�!��D���WwD�A�ڽ�*&b�������D��= (Vd���W\��V�n�U���˩n��?\]�Q�mWA[��LwYN,�96�A4��^C�� �QO� k�`�-�����'��h��aeB"�L��O�����֖g�d�����?V��Ę�ԶF}�s@���J��/kz�T9, -S^KϹC9���